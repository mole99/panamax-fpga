module manual_routing ();
endmodule
