VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO res_div
  CLASS BLOCK ;
  FOREIGN res_div ;
  ORIGIN 0.005 0.005 ;
  SIZE 56.260 BY 40.750 ;
  PIN vdda
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 0.995 36.995 3.100 39.745 ;
    END
  END vdda
  PIN vssa
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 0.995 0.995 3.100 3.745 ;
    END
  END vssa
  PIN vref
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 53.150 19.000 55.255 21.750 ;
    END
  END vref
  OBS
      LAYER pwell ;
        RECT -0.005 40.255 56.255 40.745 ;
        RECT -0.005 0.485 0.485 40.255 ;
        RECT 55.765 0.485 56.255 40.255 ;
        RECT -0.005 -0.005 56.255 0.485 ;
      LAYER li1 ;
        RECT 0.125 40.385 56.125 40.615 ;
        RECT 0.125 0.355 0.355 40.385 ;
        RECT 0.965 36.945 3.145 39.795 ;
        RECT 53.105 36.945 55.285 39.795 ;
        RECT 0.965 32.945 3.145 35.795 ;
        RECT 53.105 32.945 55.285 35.795 ;
        RECT 0.965 28.945 3.145 31.795 ;
        RECT 53.105 28.945 55.285 31.795 ;
        RECT 0.965 24.945 3.145 27.795 ;
        RECT 53.105 24.945 55.285 27.795 ;
        RECT 0.965 20.945 3.145 23.795 ;
        RECT 53.105 20.945 55.285 23.795 ;
        RECT 0.965 16.945 3.145 19.795 ;
        RECT 53.105 16.945 55.285 19.795 ;
        RECT 0.965 12.945 3.145 15.795 ;
        RECT 53.105 12.945 55.285 15.795 ;
        RECT 0.965 8.945 3.145 11.795 ;
        RECT 53.105 8.945 55.285 11.795 ;
        RECT 0.965 4.945 3.145 7.795 ;
        RECT 53.105 4.945 55.285 7.795 ;
        RECT 0.965 0.945 3.145 3.795 ;
        RECT 53.105 0.945 55.285 3.795 ;
        RECT 55.895 0.355 56.125 40.385 ;
        RECT 0.125 0.125 56.125 0.355 ;
      LAYER met1 ;
        RECT 0.125 40.385 56.125 40.615 ;
        RECT 0.125 3.745 0.355 40.385 ;
        RECT 0.995 36.995 3.100 39.745 ;
        RECT 0.995 28.995 3.100 35.745 ;
        RECT 53.150 32.995 55.255 39.745 ;
        RECT 0.995 20.995 3.100 27.745 ;
        RECT 53.150 24.995 55.255 31.745 ;
        RECT 0.995 12.995 3.100 19.745 ;
        RECT 53.150 16.995 55.255 23.745 ;
        RECT 0.995 4.995 3.100 11.745 ;
        RECT 53.150 8.995 55.255 15.745 ;
        RECT 0.125 0.355 3.100 3.745 ;
        RECT 53.150 0.995 55.255 7.745 ;
        RECT 55.895 0.355 56.125 40.385 ;
        RECT 0.125 0.125 56.125 0.355 ;
  END
END res_div
END LIBRARY

