module manual_routing (
    `ifdef USE_POWER_PINS
    inout DVPWR,
    inout DVGND
    `endif
);

endmodule
