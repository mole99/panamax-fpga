module dll (dco,
    enable,
    osc,
    resetb,
    clockp,
    div,
    ext_trim);
 input dco;
 input enable;
 input osc;
 input resetb;
 output [1:0] clockp;
 input [7:0] div;
 input [25:0] ext_trim;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire _374_;
 wire _375_;
 wire _376_;
 wire _377_;
 wire _378_;
 wire _379_;
 wire _380_;
 wire _381_;
 wire _382_;
 wire _383_;
 wire _384_;
 wire _385_;
 wire _386_;
 wire _387_;
 wire _388_;
 wire _389_;
 wire _390_;
 wire _391_;
 wire _392_;
 wire _393_;
 wire _394_;
 wire _395_;
 wire _396_;
 wire _397_;
 wire _398_;
 wire _399_;
 wire _400_;
 wire _401_;
 wire _402_;
 wire _403_;
 wire _404_;
 wire _405_;
 wire _406_;
 wire _407_;
 wire _408_;
 wire _409_;
 wire _410_;
 wire \clockp_buffer_in[0] ;
 wire \clockp_buffer_in[1] ;
 wire \dll_control.accum[0] ;
 wire \dll_control.accum[1] ;
 wire \dll_control.accum[2] ;
 wire \dll_control.accum[3] ;
 wire \dll_control.accum[4] ;
 wire \dll_control.accum[5] ;
 wire \dll_control.accum[6] ;
 wire \dll_control.accum[7] ;
 wire \dll_control.accum[8] ;
 wire \dll_control.count0[0] ;
 wire \dll_control.count0[1] ;
 wire \dll_control.count0[2] ;
 wire \dll_control.count0[3] ;
 wire \dll_control.count0[4] ;
 wire \dll_control.count0[5] ;
 wire \dll_control.count1[0] ;
 wire \dll_control.count1[1] ;
 wire \dll_control.count1[2] ;
 wire \dll_control.count1[3] ;
 wire \dll_control.count1[4] ;
 wire \dll_control.count1[5] ;
 wire \dll_control.count2[0] ;
 wire \dll_control.count2[1] ;
 wire \dll_control.count2[2] ;
 wire \dll_control.count2[3] ;
 wire \dll_control.count2[4] ;
 wire \dll_control.count2[5] ;
 wire \dll_control.count3[0] ;
 wire \dll_control.count3[1] ;
 wire \dll_control.count3[2] ;
 wire \dll_control.count3[3] ;
 wire \dll_control.count3[4] ;
 wire \dll_control.count3[5] ;
 wire \dll_control.count4[0] ;
 wire \dll_control.count4[1] ;
 wire \dll_control.count4[2] ;
 wire \dll_control.count4[3] ;
 wire \dll_control.count4[4] ;
 wire \dll_control.count4[5] ;
 wire \dll_control.count5[0] ;
 wire \dll_control.count5[1] ;
 wire \dll_control.count5[2] ;
 wire \dll_control.count5[3] ;
 wire \dll_control.count5[4] ;
 wire \dll_control.count5[5] ;
 wire \dll_control.count6[0] ;
 wire \dll_control.count6[1] ;
 wire \dll_control.count6[2] ;
 wire \dll_control.count6[3] ;
 wire \dll_control.count6[4] ;
 wire \dll_control.count6[5] ;
 wire \dll_control.count7[0] ;
 wire \dll_control.count7[1] ;
 wire \dll_control.count7[2] ;
 wire \dll_control.count7[3] ;
 wire \dll_control.count7[4] ;
 wire \dll_control.count7[5] ;
 wire \dll_control.count8[0] ;
 wire \dll_control.count8[1] ;
 wire \dll_control.count8[2] ;
 wire \dll_control.count8[3] ;
 wire \dll_control.count8[4] ;
 wire \dll_control.count8[5] ;
 wire \dll_control.oscbuf[0] ;
 wire \dll_control.oscbuf[1] ;
 wire \dll_control.oscbuf[2] ;
 wire \dll_control.tint[0] ;
 wire \dll_control.tint[1] ;
 wire \dll_control.tint[2] ;
 wire \dll_control.tint[3] ;
 wire \dll_control.tint[4] ;
 wire \dll_control.tval[0] ;
 wire \dll_control.tval[1] ;
 wire \dll_control.tval[2] ;
 wire ireset;
 wire \itrim[0] ;
 wire \itrim[10] ;
 wire \itrim[11] ;
 wire \itrim[12] ;
 wire \itrim[13] ;
 wire \itrim[14] ;
 wire \itrim[15] ;
 wire \itrim[16] ;
 wire \itrim[17] ;
 wire \itrim[18] ;
 wire \itrim[19] ;
 wire \itrim[1] ;
 wire \itrim[20] ;
 wire \itrim[21] ;
 wire \itrim[22] ;
 wire \itrim[23] ;
 wire \itrim[24] ;
 wire \itrim[25] ;
 wire \itrim[2] ;
 wire \itrim[3] ;
 wire \itrim[4] ;
 wire \itrim[5] ;
 wire \itrim[6] ;
 wire \itrim[7] ;
 wire \itrim[8] ;
 wire \itrim[9] ;
 wire \ringosc.c[0] ;
 wire \ringosc.c[1] ;
 wire \ringosc.dstage[0].id.d0 ;
 wire \ringosc.dstage[0].id.d1 ;
 wire \ringosc.dstage[0].id.d2 ;
 wire \ringosc.dstage[0].id.in ;
 wire \ringosc.dstage[0].id.out ;
 wire \ringosc.dstage[0].id.ts ;
 wire \ringosc.dstage[10].id.d0 ;
 wire \ringosc.dstage[10].id.d1 ;
 wire \ringosc.dstage[10].id.d2 ;
 wire \ringosc.dstage[10].id.in ;
 wire \ringosc.dstage[10].id.out ;
 wire \ringosc.dstage[10].id.ts ;
 wire \ringosc.dstage[11].id.d0 ;
 wire \ringosc.dstage[11].id.d1 ;
 wire \ringosc.dstage[11].id.d2 ;
 wire \ringosc.dstage[11].id.out ;
 wire \ringosc.dstage[11].id.ts ;
 wire \ringosc.dstage[1].id.d0 ;
 wire \ringosc.dstage[1].id.d1 ;
 wire \ringosc.dstage[1].id.d2 ;
 wire \ringosc.dstage[1].id.out ;
 wire \ringosc.dstage[1].id.ts ;
 wire \ringosc.dstage[2].id.d0 ;
 wire \ringosc.dstage[2].id.d1 ;
 wire \ringosc.dstage[2].id.d2 ;
 wire \ringosc.dstage[2].id.out ;
 wire \ringosc.dstage[2].id.ts ;
 wire \ringosc.dstage[3].id.d0 ;
 wire \ringosc.dstage[3].id.d1 ;
 wire \ringosc.dstage[3].id.d2 ;
 wire \ringosc.dstage[3].id.out ;
 wire \ringosc.dstage[3].id.ts ;
 wire \ringosc.dstage[4].id.d0 ;
 wire \ringosc.dstage[4].id.d1 ;
 wire \ringosc.dstage[4].id.d2 ;
 wire \ringosc.dstage[4].id.out ;
 wire \ringosc.dstage[4].id.ts ;
 wire \ringosc.dstage[5].id.d0 ;
 wire \ringosc.dstage[5].id.d1 ;
 wire \ringosc.dstage[5].id.d2 ;
 wire \ringosc.dstage[5].id.out ;
 wire \ringosc.dstage[5].id.ts ;
 wire \ringosc.dstage[6].id.d0 ;
 wire \ringosc.dstage[6].id.d1 ;
 wire \ringosc.dstage[6].id.d2 ;
 wire \ringosc.dstage[6].id.out ;
 wire \ringosc.dstage[6].id.ts ;
 wire \ringosc.dstage[7].id.d0 ;
 wire \ringosc.dstage[7].id.d1 ;
 wire \ringosc.dstage[7].id.d2 ;
 wire \ringosc.dstage[7].id.out ;
 wire \ringosc.dstage[7].id.ts ;
 wire \ringosc.dstage[8].id.d0 ;
 wire \ringosc.dstage[8].id.d1 ;
 wire \ringosc.dstage[8].id.d2 ;
 wire \ringosc.dstage[8].id.out ;
 wire \ringosc.dstage[8].id.ts ;
 wire \ringosc.dstage[9].id.d0 ;
 wire \ringosc.dstage[9].id.d1 ;
 wire \ringosc.dstage[9].id.d2 ;
 wire \ringosc.dstage[9].id.ts ;
 wire \ringosc.iss.ctrl0 ;
 wire \ringosc.iss.d0 ;
 wire \ringosc.iss.d1 ;
 wire \ringosc.iss.d2 ;
 wire \ringosc.iss.one ;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;

 sky130_fd_sc_hd__nand2b_1 _411_ (.A_N(\dll_control.accum[6] ),
    .B(\dll_control.accum[7] ),
    .Y(_145_));
 sky130_fd_sc_hd__nand2b_1 _412_ (.A_N(\dll_control.count8[5] ),
    .B(\dll_control.accum[5] ),
    .Y(_146_));
 sky130_fd_sc_hd__xnor2_1 _413_ (.A(\dll_control.accum[5] ),
    .B(\dll_control.count8[5] ),
    .Y(_147_));
 sky130_fd_sc_hd__nand2_1 _414_ (.A(\dll_control.count0[5] ),
    .B(_147_),
    .Y(_148_));
 sky130_fd_sc_hd__a21o_1 _415_ (.A1(_146_),
    .A2(_148_),
    .B1(\dll_control.accum[6] ),
    .X(_149_));
 sky130_fd_sc_hd__nand3_1 _416_ (.A(\dll_control.accum[6] ),
    .B(_146_),
    .C(_148_),
    .Y(_150_));
 sky130_fd_sc_hd__nand2_1 _417_ (.A(_149_),
    .B(_150_),
    .Y(_151_));
 sky130_fd_sc_hd__xnor2_1 _418_ (.A(\dll_control.count0[5] ),
    .B(_147_),
    .Y(_152_));
 sky130_fd_sc_hd__nand2b_1 _419_ (.A_N(\dll_control.count8[4] ),
    .B(\dll_control.accum[4] ),
    .Y(_153_));
 sky130_fd_sc_hd__xnor2_1 _420_ (.A(\dll_control.accum[4] ),
    .B(\dll_control.count8[4] ),
    .Y(_154_));
 sky130_fd_sc_hd__nand2_1 _421_ (.A(\dll_control.count0[4] ),
    .B(_154_),
    .Y(_155_));
 sky130_fd_sc_hd__nand3_1 _422_ (.A(_152_),
    .B(_153_),
    .C(_155_),
    .Y(_156_));
 sky130_fd_sc_hd__xnor2_1 _423_ (.A(\dll_control.accum[3] ),
    .B(\dll_control.count8[3] ),
    .Y(_157_));
 sky130_fd_sc_hd__xnor2_1 _424_ (.A(\dll_control.count0[3] ),
    .B(_157_),
    .Y(_158_));
 sky130_fd_sc_hd__nand2b_1 _425_ (.A_N(\dll_control.count8[2] ),
    .B(\dll_control.accum[2] ),
    .Y(_159_));
 sky130_fd_sc_hd__xnor2_1 _426_ (.A(\dll_control.accum[2] ),
    .B(\dll_control.count8[2] ),
    .Y(_160_));
 sky130_fd_sc_hd__nand2_1 _427_ (.A(\dll_control.count0[2] ),
    .B(_160_),
    .Y(_161_));
 sky130_fd_sc_hd__nand3_1 _428_ (.A(_158_),
    .B(_159_),
    .C(_161_),
    .Y(_162_));
 sky130_fd_sc_hd__xor2_1 _429_ (.A(\dll_control.count8[0] ),
    .B(\dll_control.count0[0] ),
    .X(_163_));
 sky130_fd_sc_hd__and2b_1 _430_ (.A_N(\dll_control.count0[0] ),
    .B(\dll_control.count8[0] ),
    .X(_164_));
 sky130_fd_sc_hd__xnor2_1 _431_ (.A(\dll_control.accum[1] ),
    .B(\dll_control.count8[1] ),
    .Y(_165_));
 sky130_fd_sc_hd__xnor2_1 _432_ (.A(\dll_control.count0[1] ),
    .B(_165_),
    .Y(_166_));
 sky130_fd_sc_hd__xor2_1 _433_ (.A(_164_),
    .B(_166_),
    .X(_167_));
 sky130_fd_sc_hd__nor2_1 _434_ (.A(_164_),
    .B(_166_),
    .Y(_168_));
 sky130_fd_sc_hd__a31o_1 _435_ (.A1(\dll_control.accum[0] ),
    .A2(_163_),
    .A3(_167_),
    .B1(_168_),
    .X(_169_));
 sky130_fd_sc_hd__xnor2_1 _436_ (.A(\dll_control.count0[2] ),
    .B(_160_),
    .Y(_170_));
 sky130_fd_sc_hd__nand2b_1 _437_ (.A_N(\dll_control.count8[1] ),
    .B(\dll_control.accum[1] ),
    .Y(_171_));
 sky130_fd_sc_hd__nand2_1 _438_ (.A(\dll_control.count0[1] ),
    .B(_165_),
    .Y(_172_));
 sky130_fd_sc_hd__nand3_1 _439_ (.A(_170_),
    .B(_171_),
    .C(_172_),
    .Y(_173_));
 sky130_fd_sc_hd__a21oi_1 _440_ (.A1(_171_),
    .A2(_172_),
    .B1(_170_),
    .Y(_174_));
 sky130_fd_sc_hd__a21o_1 _441_ (.A1(_169_),
    .A2(_173_),
    .B1(_174_),
    .X(_175_));
 sky130_fd_sc_hd__a21oi_1 _442_ (.A1(_159_),
    .A2(_161_),
    .B1(_158_),
    .Y(_176_));
 sky130_fd_sc_hd__a21oi_1 _443_ (.A1(_162_),
    .A2(_175_),
    .B1(_176_),
    .Y(_177_));
 sky130_fd_sc_hd__nand2b_1 _444_ (.A_N(\dll_control.count8[3] ),
    .B(\dll_control.accum[3] ),
    .Y(_178_));
 sky130_fd_sc_hd__nand2_1 _445_ (.A(\dll_control.count0[3] ),
    .B(_157_),
    .Y(_179_));
 sky130_fd_sc_hd__xnor2_1 _446_ (.A(\dll_control.count0[4] ),
    .B(_154_),
    .Y(_180_));
 sky130_fd_sc_hd__a21o_1 _447_ (.A1(_178_),
    .A2(_179_),
    .B1(_180_),
    .X(_181_));
 sky130_fd_sc_hd__nand3_1 _448_ (.A(_180_),
    .B(_178_),
    .C(_179_),
    .Y(_182_));
 sky130_fd_sc_hd__nand2_1 _449_ (.A(_181_),
    .B(_182_),
    .Y(_183_));
 sky130_fd_sc_hd__o21ai_1 _450_ (.A1(_177_),
    .A2(_183_),
    .B1(_181_),
    .Y(_184_));
 sky130_fd_sc_hd__a21oi_1 _451_ (.A1(_153_),
    .A2(_155_),
    .B1(_152_),
    .Y(_185_));
 sky130_fd_sc_hd__a21oi_1 _452_ (.A1(_156_),
    .A2(_184_),
    .B1(_185_),
    .Y(_186_));
 sky130_fd_sc_hd__o21ai_1 _453_ (.A1(_151_),
    .A2(_186_),
    .B1(_149_),
    .Y(_187_));
 sky130_fd_sc_hd__and2b_1 _454_ (.A_N(\dll_control.accum[7] ),
    .B(\dll_control.accum[6] ),
    .X(_188_));
 sky130_fd_sc_hd__a21oi_1 _455_ (.A1(_145_),
    .A2(_187_),
    .B1(_188_),
    .Y(_189_));
 sky130_fd_sc_hd__xnor2_1 _456_ (.A(\dll_control.accum[8] ),
    .B(\dll_control.accum[7] ),
    .Y(_190_));
 sky130_fd_sc_hd__xnor2_1 _457_ (.A(_189_),
    .B(_190_),
    .Y(_191_));
 sky130_fd_sc_hd__and2b_1 _458_ (.A_N(\dll_control.oscbuf[1] ),
    .B(\dll_control.oscbuf[2] ),
    .X(_192_));
 sky130_fd_sc_hd__clkbuf_2 _459_ (.A(_192_),
    .X(_193_));
 sky130_fd_sc_hd__buf_2 _460_ (.A(_193_),
    .X(_194_));
 sky130_fd_sc_hd__mux2_1 _461_ (.A0(\dll_control.accum[8] ),
    .A1(_191_),
    .S(_194_),
    .X(_195_));
 sky130_fd_sc_hd__clkbuf_1 _462_ (.A(_195_),
    .X(_144_));
 sky130_fd_sc_hd__nand2b_1 _463_ (.A_N(_188_),
    .B(_145_),
    .Y(_196_));
 sky130_fd_sc_hd__xnor2_1 _464_ (.A(_196_),
    .B(_187_),
    .Y(_197_));
 sky130_fd_sc_hd__mux2_1 _465_ (.A0(\dll_control.accum[7] ),
    .A1(_197_),
    .S(_194_),
    .X(_198_));
 sky130_fd_sc_hd__clkbuf_1 _466_ (.A(_198_),
    .X(_143_));
 sky130_fd_sc_hd__xor2_1 _467_ (.A(_151_),
    .B(_186_),
    .X(_199_));
 sky130_fd_sc_hd__mux2_1 _468_ (.A0(\dll_control.accum[6] ),
    .A1(_199_),
    .S(_194_),
    .X(_200_));
 sky130_fd_sc_hd__clkbuf_1 _469_ (.A(_200_),
    .X(_142_));
 sky130_fd_sc_hd__nand2b_1 _470_ (.A_N(_185_),
    .B(_156_),
    .Y(_201_));
 sky130_fd_sc_hd__xnor2_1 _471_ (.A(_201_),
    .B(_184_),
    .Y(_202_));
 sky130_fd_sc_hd__mux2_1 _472_ (.A0(\dll_control.accum[5] ),
    .A1(_202_),
    .S(_194_),
    .X(_203_));
 sky130_fd_sc_hd__clkbuf_1 _473_ (.A(_203_),
    .X(_141_));
 sky130_fd_sc_hd__xor2_1 _474_ (.A(_177_),
    .B(_183_),
    .X(_204_));
 sky130_fd_sc_hd__mux2_1 _475_ (.A0(\dll_control.accum[4] ),
    .A1(_204_),
    .S(_194_),
    .X(_205_));
 sky130_fd_sc_hd__clkbuf_1 _476_ (.A(_205_),
    .X(_140_));
 sky130_fd_sc_hd__nand2b_1 _477_ (.A_N(_176_),
    .B(_162_),
    .Y(_206_));
 sky130_fd_sc_hd__xnor2_1 _478_ (.A(_206_),
    .B(_175_),
    .Y(_207_));
 sky130_fd_sc_hd__mux2_1 _479_ (.A0(\dll_control.accum[3] ),
    .A1(_207_),
    .S(_194_),
    .X(_208_));
 sky130_fd_sc_hd__clkbuf_1 _480_ (.A(_208_),
    .X(_139_));
 sky130_fd_sc_hd__nand2b_1 _481_ (.A_N(_174_),
    .B(_173_),
    .Y(_209_));
 sky130_fd_sc_hd__xnor2_1 _482_ (.A(_169_),
    .B(_209_),
    .Y(_210_));
 sky130_fd_sc_hd__buf_2 _483_ (.A(_193_),
    .X(_211_));
 sky130_fd_sc_hd__mux2_1 _484_ (.A0(\dll_control.accum[2] ),
    .A1(_210_),
    .S(_211_),
    .X(_212_));
 sky130_fd_sc_hd__clkbuf_1 _485_ (.A(_212_),
    .X(_138_));
 sky130_fd_sc_hd__nand2_1 _486_ (.A(\dll_control.accum[0] ),
    .B(_163_),
    .Y(_213_));
 sky130_fd_sc_hd__xnor2_1 _487_ (.A(_213_),
    .B(_167_),
    .Y(_214_));
 sky130_fd_sc_hd__mux2_1 _488_ (.A0(\dll_control.accum[1] ),
    .A1(_214_),
    .S(_211_),
    .X(_215_));
 sky130_fd_sc_hd__clkbuf_1 _489_ (.A(_215_),
    .X(_137_));
 sky130_fd_sc_hd__nand2b_1 _490_ (.A_N(\dll_control.oscbuf[1] ),
    .B(\dll_control.oscbuf[2] ),
    .Y(_216_));
 sky130_fd_sc_hd__buf_2 _491_ (.A(_216_),
    .X(_217_));
 sky130_fd_sc_hd__clkbuf_2 _492_ (.A(_217_),
    .X(_218_));
 sky130_fd_sc_hd__a21o_1 _493_ (.A1(_194_),
    .A2(_163_),
    .B1(\dll_control.accum[0] ),
    .X(_219_));
 sky130_fd_sc_hd__o21a_1 _494_ (.A1(_218_),
    .A2(_213_),
    .B1(_219_),
    .X(_136_));
 sky130_fd_sc_hd__mux2_1 _495_ (.A0(\dll_control.count4[5] ),
    .A1(\dll_control.count3[5] ),
    .S(_211_),
    .X(_220_));
 sky130_fd_sc_hd__clkbuf_1 _496_ (.A(_220_),
    .X(_135_));
 sky130_fd_sc_hd__mux2_1 _497_ (.A0(\dll_control.count4[4] ),
    .A1(\dll_control.count3[4] ),
    .S(_211_),
    .X(_221_));
 sky130_fd_sc_hd__clkbuf_1 _498_ (.A(_221_),
    .X(_134_));
 sky130_fd_sc_hd__mux2_1 _499_ (.A0(\dll_control.count4[3] ),
    .A1(\dll_control.count3[3] ),
    .S(_211_),
    .X(_222_));
 sky130_fd_sc_hd__clkbuf_1 _500_ (.A(_222_),
    .X(_133_));
 sky130_fd_sc_hd__mux2_1 _501_ (.A0(\dll_control.count4[2] ),
    .A1(\dll_control.count3[2] ),
    .S(_211_),
    .X(_223_));
 sky130_fd_sc_hd__clkbuf_1 _502_ (.A(_223_),
    .X(_132_));
 sky130_fd_sc_hd__mux2_1 _503_ (.A0(\dll_control.count4[1] ),
    .A1(\dll_control.count3[1] ),
    .S(_211_),
    .X(_224_));
 sky130_fd_sc_hd__clkbuf_1 _504_ (.A(_224_),
    .X(_131_));
 sky130_fd_sc_hd__buf_2 _505_ (.A(_193_),
    .X(_225_));
 sky130_fd_sc_hd__mux2_1 _506_ (.A0(\dll_control.count4[0] ),
    .A1(\dll_control.count3[0] ),
    .S(_225_),
    .X(_226_));
 sky130_fd_sc_hd__clkbuf_1 _507_ (.A(_226_),
    .X(_130_));
 sky130_fd_sc_hd__mux2_1 _508_ (.A0(\dll_control.count8[5] ),
    .A1(\dll_control.count7[5] ),
    .S(_225_),
    .X(_227_));
 sky130_fd_sc_hd__clkbuf_1 _509_ (.A(_227_),
    .X(_129_));
 sky130_fd_sc_hd__mux2_1 _510_ (.A0(\dll_control.count8[4] ),
    .A1(\dll_control.count7[4] ),
    .S(_225_),
    .X(_228_));
 sky130_fd_sc_hd__clkbuf_1 _511_ (.A(_228_),
    .X(_128_));
 sky130_fd_sc_hd__mux2_1 _512_ (.A0(\dll_control.count8[3] ),
    .A1(\dll_control.count7[3] ),
    .S(_225_),
    .X(_229_));
 sky130_fd_sc_hd__clkbuf_1 _513_ (.A(_229_),
    .X(_127_));
 sky130_fd_sc_hd__mux2_1 _514_ (.A0(\dll_control.count8[2] ),
    .A1(\dll_control.count7[2] ),
    .S(_225_),
    .X(_230_));
 sky130_fd_sc_hd__clkbuf_1 _515_ (.A(_230_),
    .X(_126_));
 sky130_fd_sc_hd__mux2_1 _516_ (.A0(\dll_control.count8[1] ),
    .A1(\dll_control.count7[1] ),
    .S(_225_),
    .X(_231_));
 sky130_fd_sc_hd__clkbuf_1 _517_ (.A(_231_),
    .X(_125_));
 sky130_fd_sc_hd__mux2_1 _518_ (.A0(\dll_control.count8[0] ),
    .A1(\dll_control.count7[0] ),
    .S(_225_),
    .X(_232_));
 sky130_fd_sc_hd__clkbuf_1 _519_ (.A(_232_),
    .X(_124_));
 sky130_fd_sc_hd__buf_2 _520_ (.A(_193_),
    .X(_233_));
 sky130_fd_sc_hd__mux2_1 _521_ (.A0(\dll_control.count3[5] ),
    .A1(\dll_control.count2[5] ),
    .S(_233_),
    .X(_234_));
 sky130_fd_sc_hd__clkbuf_1 _522_ (.A(_234_),
    .X(_123_));
 sky130_fd_sc_hd__mux2_1 _523_ (.A0(\dll_control.count3[4] ),
    .A1(\dll_control.count2[4] ),
    .S(_233_),
    .X(_235_));
 sky130_fd_sc_hd__clkbuf_1 _524_ (.A(_235_),
    .X(_122_));
 sky130_fd_sc_hd__mux2_1 _525_ (.A0(\dll_control.count3[3] ),
    .A1(\dll_control.count2[3] ),
    .S(_233_),
    .X(_236_));
 sky130_fd_sc_hd__clkbuf_1 _526_ (.A(_236_),
    .X(_121_));
 sky130_fd_sc_hd__mux2_1 _527_ (.A0(\dll_control.count3[2] ),
    .A1(\dll_control.count2[2] ),
    .S(_233_),
    .X(_237_));
 sky130_fd_sc_hd__clkbuf_1 _528_ (.A(_237_),
    .X(_120_));
 sky130_fd_sc_hd__mux2_1 _529_ (.A0(\dll_control.count3[1] ),
    .A1(\dll_control.count2[1] ),
    .S(_233_),
    .X(_238_));
 sky130_fd_sc_hd__clkbuf_1 _530_ (.A(_238_),
    .X(_119_));
 sky130_fd_sc_hd__mux2_1 _531_ (.A0(\dll_control.count3[0] ),
    .A1(\dll_control.count2[0] ),
    .S(_233_),
    .X(_239_));
 sky130_fd_sc_hd__clkbuf_1 _532_ (.A(_239_),
    .X(_118_));
 sky130_fd_sc_hd__mux2_1 _533_ (.A0(\dll_control.count7[5] ),
    .A1(\dll_control.count6[5] ),
    .S(_233_),
    .X(_240_));
 sky130_fd_sc_hd__clkbuf_1 _534_ (.A(_240_),
    .X(_117_));
 sky130_fd_sc_hd__buf_2 _535_ (.A(_192_),
    .X(_241_));
 sky130_fd_sc_hd__mux2_1 _536_ (.A0(\dll_control.count7[4] ),
    .A1(\dll_control.count6[4] ),
    .S(_241_),
    .X(_242_));
 sky130_fd_sc_hd__clkbuf_1 _537_ (.A(_242_),
    .X(_116_));
 sky130_fd_sc_hd__mux2_1 _538_ (.A0(\dll_control.count7[3] ),
    .A1(\dll_control.count6[3] ),
    .S(_241_),
    .X(_243_));
 sky130_fd_sc_hd__clkbuf_1 _539_ (.A(_243_),
    .X(_115_));
 sky130_fd_sc_hd__mux2_1 _540_ (.A0(\dll_control.count7[2] ),
    .A1(\dll_control.count6[2] ),
    .S(_241_),
    .X(_244_));
 sky130_fd_sc_hd__clkbuf_1 _541_ (.A(_244_),
    .X(_114_));
 sky130_fd_sc_hd__mux2_1 _542_ (.A0(\dll_control.count7[1] ),
    .A1(\dll_control.count6[1] ),
    .S(_241_),
    .X(_245_));
 sky130_fd_sc_hd__clkbuf_1 _543_ (.A(_245_),
    .X(_113_));
 sky130_fd_sc_hd__mux2_1 _544_ (.A0(\dll_control.count7[0] ),
    .A1(\dll_control.count6[0] ),
    .S(_241_),
    .X(_246_));
 sky130_fd_sc_hd__clkbuf_1 _545_ (.A(_246_),
    .X(_112_));
 sky130_fd_sc_hd__and3_1 _546_ (.A(\dll_control.count0[2] ),
    .B(\dll_control.count0[1] ),
    .C(\dll_control.count0[0] ),
    .X(_247_));
 sky130_fd_sc_hd__and3_1 _547_ (.A(\dll_control.count0[4] ),
    .B(\dll_control.count0[3] ),
    .C(_247_),
    .X(_248_));
 sky130_fd_sc_hd__o21a_1 _548_ (.A1(\dll_control.count0[5] ),
    .A2(_248_),
    .B1(_218_),
    .X(_111_));
 sky130_fd_sc_hd__inv_1 _549_ (.A(_248_),
    .Y(_249_));
 sky130_fd_sc_hd__a21o_1 _550_ (.A1(\dll_control.count0[3] ),
    .A2(_247_),
    .B1(\dll_control.count0[4] ),
    .X(_250_));
 sky130_fd_sc_hd__o211a_1 _551_ (.A1(\dll_control.count0[5] ),
    .A2(_249_),
    .B1(_250_),
    .C1(_218_),
    .X(_110_));
 sky130_fd_sc_hd__xor2_1 _552_ (.A(\dll_control.count0[3] ),
    .B(_247_),
    .X(_251_));
 sky130_fd_sc_hd__clkbuf_2 _553_ (.A(_216_),
    .X(_252_));
 sky130_fd_sc_hd__and3_1 _554_ (.A(\dll_control.count0[5] ),
    .B(_252_),
    .C(_248_),
    .X(_253_));
 sky130_fd_sc_hd__a21o_1 _555_ (.A1(_218_),
    .A2(_251_),
    .B1(_253_),
    .X(_109_));
 sky130_fd_sc_hd__a21oi_1 _556_ (.A1(\dll_control.count0[1] ),
    .A2(\dll_control.count0[0] ),
    .B1(\dll_control.count0[2] ),
    .Y(_254_));
 sky130_fd_sc_hd__nor2_1 _557_ (.A(_247_),
    .B(_254_),
    .Y(_255_));
 sky130_fd_sc_hd__a21o_1 _558_ (.A1(_218_),
    .A2(_255_),
    .B1(_253_),
    .X(_108_));
 sky130_fd_sc_hd__xor2_1 _559_ (.A(\dll_control.count0[1] ),
    .B(\dll_control.count0[0] ),
    .X(_256_));
 sky130_fd_sc_hd__a21o_1 _560_ (.A1(_218_),
    .A2(_256_),
    .B1(_253_),
    .X(_107_));
 sky130_fd_sc_hd__nand3b_1 _561_ (.A_N(_253_),
    .B(\dll_control.count0[0] ),
    .C(_218_),
    .Y(_106_));
 sky130_fd_sc_hd__mux2_1 _562_ (.A0(\dll_control.count4[5] ),
    .A1(\dll_control.count5[5] ),
    .S(_217_),
    .X(_257_));
 sky130_fd_sc_hd__clkbuf_1 _563_ (.A(_257_),
    .X(_105_));
 sky130_fd_sc_hd__mux2_1 _564_ (.A0(\dll_control.count4[4] ),
    .A1(\dll_control.count5[4] ),
    .S(_217_),
    .X(_258_));
 sky130_fd_sc_hd__clkbuf_1 _565_ (.A(_258_),
    .X(_104_));
 sky130_fd_sc_hd__mux2_1 _566_ (.A0(\dll_control.count4[3] ),
    .A1(\dll_control.count5[3] ),
    .S(_217_),
    .X(_259_));
 sky130_fd_sc_hd__clkbuf_1 _567_ (.A(_259_),
    .X(_103_));
 sky130_fd_sc_hd__mux2_1 _568_ (.A0(\dll_control.count4[2] ),
    .A1(\dll_control.count5[2] ),
    .S(_217_),
    .X(_260_));
 sky130_fd_sc_hd__clkbuf_1 _569_ (.A(_260_),
    .X(_102_));
 sky130_fd_sc_hd__mux2_1 _570_ (.A0(\dll_control.count4[1] ),
    .A1(\dll_control.count5[1] ),
    .S(_217_),
    .X(_261_));
 sky130_fd_sc_hd__clkbuf_1 _571_ (.A(_261_),
    .X(_101_));
 sky130_fd_sc_hd__mux2_1 _572_ (.A0(\dll_control.count4[0] ),
    .A1(\dll_control.count5[0] ),
    .S(_217_),
    .X(_262_));
 sky130_fd_sc_hd__clkbuf_1 _573_ (.A(_262_),
    .X(_100_));
 sky130_fd_sc_hd__mux2_1 _574_ (.A0(\dll_control.count0[5] ),
    .A1(\dll_control.count1[5] ),
    .S(_252_),
    .X(_263_));
 sky130_fd_sc_hd__clkbuf_1 _575_ (.A(_263_),
    .X(_099_));
 sky130_fd_sc_hd__mux2_1 _576_ (.A0(\dll_control.count0[4] ),
    .A1(\dll_control.count1[4] ),
    .S(_252_),
    .X(_264_));
 sky130_fd_sc_hd__clkbuf_1 _577_ (.A(_264_),
    .X(_098_));
 sky130_fd_sc_hd__mux2_1 _578_ (.A0(\dll_control.count0[3] ),
    .A1(\dll_control.count1[3] ),
    .S(_252_),
    .X(_265_));
 sky130_fd_sc_hd__clkbuf_1 _579_ (.A(_265_),
    .X(_097_));
 sky130_fd_sc_hd__mux2_1 _580_ (.A0(\dll_control.count0[2] ),
    .A1(\dll_control.count1[2] ),
    .S(_252_),
    .X(_266_));
 sky130_fd_sc_hd__clkbuf_1 _581_ (.A(_266_),
    .X(_096_));
 sky130_fd_sc_hd__mux2_1 _582_ (.A0(\dll_control.count0[1] ),
    .A1(\dll_control.count1[1] ),
    .S(_252_),
    .X(_267_));
 sky130_fd_sc_hd__clkbuf_1 _583_ (.A(_267_),
    .X(_095_));
 sky130_fd_sc_hd__mux2_1 _584_ (.A0(\dll_control.count0[0] ),
    .A1(\dll_control.count1[0] ),
    .S(_252_),
    .X(_268_));
 sky130_fd_sc_hd__clkbuf_1 _585_ (.A(_268_),
    .X(_094_));
 sky130_fd_sc_hd__mux2_1 _586_ (.A0(\dll_control.count6[5] ),
    .A1(\dll_control.count5[5] ),
    .S(_241_),
    .X(_269_));
 sky130_fd_sc_hd__clkbuf_1 _587_ (.A(_269_),
    .X(_093_));
 sky130_fd_sc_hd__mux2_1 _588_ (.A0(\dll_control.count6[4] ),
    .A1(\dll_control.count5[4] ),
    .S(_241_),
    .X(_270_));
 sky130_fd_sc_hd__clkbuf_1 _589_ (.A(_270_),
    .X(_092_));
 sky130_fd_sc_hd__buf_2 _590_ (.A(_192_),
    .X(_271_));
 sky130_fd_sc_hd__mux2_1 _591_ (.A0(\dll_control.count6[3] ),
    .A1(\dll_control.count5[3] ),
    .S(_271_),
    .X(_272_));
 sky130_fd_sc_hd__clkbuf_1 _592_ (.A(_272_),
    .X(_091_));
 sky130_fd_sc_hd__mux2_1 _593_ (.A0(\dll_control.count6[2] ),
    .A1(\dll_control.count5[2] ),
    .S(_271_),
    .X(_273_));
 sky130_fd_sc_hd__clkbuf_1 _594_ (.A(_273_),
    .X(_090_));
 sky130_fd_sc_hd__mux2_1 _595_ (.A0(\dll_control.count6[1] ),
    .A1(\dll_control.count5[1] ),
    .S(_271_),
    .X(_274_));
 sky130_fd_sc_hd__clkbuf_1 _596_ (.A(_274_),
    .X(_089_));
 sky130_fd_sc_hd__mux2_1 _597_ (.A0(\dll_control.count6[0] ),
    .A1(\dll_control.count5[0] ),
    .S(_271_),
    .X(_275_));
 sky130_fd_sc_hd__clkbuf_1 _598_ (.A(_275_),
    .X(_088_));
 sky130_fd_sc_hd__mux2_1 _599_ (.A0(\dll_control.count2[5] ),
    .A1(\dll_control.count1[5] ),
    .S(_271_),
    .X(_276_));
 sky130_fd_sc_hd__clkbuf_1 _600_ (.A(_276_),
    .X(_087_));
 sky130_fd_sc_hd__mux2_1 _601_ (.A0(\dll_control.count2[4] ),
    .A1(\dll_control.count1[4] ),
    .S(_271_),
    .X(_277_));
 sky130_fd_sc_hd__clkbuf_1 _602_ (.A(_277_),
    .X(_086_));
 sky130_fd_sc_hd__mux2_1 _603_ (.A0(\dll_control.count2[3] ),
    .A1(\dll_control.count1[3] ),
    .S(_271_),
    .X(_278_));
 sky130_fd_sc_hd__clkbuf_1 _604_ (.A(_278_),
    .X(_085_));
 sky130_fd_sc_hd__mux2_1 _605_ (.A0(\dll_control.count2[2] ),
    .A1(\dll_control.count1[2] ),
    .S(_193_),
    .X(_279_));
 sky130_fd_sc_hd__clkbuf_1 _606_ (.A(_279_),
    .X(_084_));
 sky130_fd_sc_hd__mux2_1 _607_ (.A0(\dll_control.count2[1] ),
    .A1(\dll_control.count1[1] ),
    .S(_193_),
    .X(_280_));
 sky130_fd_sc_hd__clkbuf_1 _608_ (.A(_280_),
    .X(_083_));
 sky130_fd_sc_hd__mux2_1 _609_ (.A0(\dll_control.count2[0] ),
    .A1(\dll_control.count1[0] ),
    .S(_193_),
    .X(_281_));
 sky130_fd_sc_hd__clkbuf_1 _610_ (.A(_281_),
    .X(_082_));
 sky130_fd_sc_hd__inv_2 _611_ (.A(div[5]),
    .Y(_282_));
 sky130_fd_sc_hd__inv_2 _612_ (.A(div[4]),
    .Y(_283_));
 sky130_fd_sc_hd__o22a_1 _613_ (.A1(\dll_control.accum[5] ),
    .A2(_282_),
    .B1(_283_),
    .B2(\dll_control.accum[4] ),
    .X(_284_));
 sky130_fd_sc_hd__and2_1 _614_ (.A(\dll_control.accum[5] ),
    .B(_282_),
    .X(_285_));
 sky130_fd_sc_hd__nand2b_1 _615_ (.A_N(\dll_control.accum[6] ),
    .B(div[6]),
    .Y(_286_));
 sky130_fd_sc_hd__nand2b_1 _616_ (.A_N(\dll_control.accum[7] ),
    .B(div[7]),
    .Y(_287_));
 sky130_fd_sc_hd__nand2b_1 _617_ (.A_N(div[7]),
    .B(\dll_control.accum[7] ),
    .Y(_288_));
 sky130_fd_sc_hd__nand2b_1 _618_ (.A_N(div[6]),
    .B(\dll_control.accum[6] ),
    .Y(_289_));
 sky130_fd_sc_hd__nand4_1 _619_ (.A(_286_),
    .B(_287_),
    .C(_288_),
    .D(_289_),
    .Y(_290_));
 sky130_fd_sc_hd__and2b_1 _620_ (.A_N(div[7]),
    .B(\dll_control.accum[7] ),
    .X(_291_));
 sky130_fd_sc_hd__o21a_1 _621_ (.A1(_286_),
    .A2(_291_),
    .B1(_287_),
    .X(_292_));
 sky130_fd_sc_hd__o31a_1 _622_ (.A1(_284_),
    .A2(_285_),
    .A3(_290_),
    .B1(_292_),
    .X(_293_));
 sky130_fd_sc_hd__a21oi_1 _623_ (.A1(\dll_control.accum[4] ),
    .A2(_283_),
    .B1(\dll_control.accum[8] ),
    .Y(_294_));
 sky130_fd_sc_hd__and4bb_1 _624_ (.A_N(_285_),
    .B_N(_290_),
    .C(_294_),
    .D(_284_),
    .X(_295_));
 sky130_fd_sc_hd__inv_1 _625_ (.A(\dll_control.accum[3] ),
    .Y(_296_));
 sky130_fd_sc_hd__nand2b_1 _626_ (.A_N(\dll_control.accum[3] ),
    .B(div[3]),
    .Y(_297_));
 sky130_fd_sc_hd__nand2b_1 _627_ (.A_N(div[3]),
    .B(\dll_control.accum[3] ),
    .Y(_298_));
 sky130_fd_sc_hd__xnor2_1 _628_ (.A(\dll_control.accum[2] ),
    .B(div[2]),
    .Y(_299_));
 sky130_fd_sc_hd__and3_1 _629_ (.A(_297_),
    .B(_298_),
    .C(_299_),
    .X(_300_));
 sky130_fd_sc_hd__nand2b_1 _630_ (.A_N(div[0]),
    .B(\dll_control.accum[0] ),
    .Y(_301_));
 sky130_fd_sc_hd__nand2b_1 _631_ (.A_N(div[1]),
    .B(\dll_control.accum[1] ),
    .Y(_302_));
 sky130_fd_sc_hd__and2b_1 _632_ (.A_N(\dll_control.accum[1] ),
    .B(div[1]),
    .X(_303_));
 sky130_fd_sc_hd__a21o_1 _633_ (.A1(_301_),
    .A2(_302_),
    .B1(_303_),
    .X(_304_));
 sky130_fd_sc_hd__and3b_1 _634_ (.A_N(\dll_control.accum[2] ),
    .B(div[2]),
    .C(_298_),
    .X(_305_));
 sky130_fd_sc_hd__a221o_1 _635_ (.A1(_296_),
    .A2(div[3]),
    .B1(_300_),
    .B2(_304_),
    .C1(_305_),
    .X(_306_));
 sky130_fd_sc_hd__a2bb2o_2 _636_ (.A1_N(\dll_control.accum[8] ),
    .A2_N(_293_),
    .B1(_295_),
    .B2(_306_),
    .X(_307_));
 sky130_fd_sc_hd__clkbuf_2 _637_ (.A(_307_),
    .X(_308_));
 sky130_fd_sc_hd__nor2_1 _638_ (.A(net110),
    .B(_308_),
    .Y(_309_));
 sky130_fd_sc_hd__nor2_1 _639_ (.A(net111),
    .B(_308_),
    .Y(_310_));
 sky130_fd_sc_hd__nor2_1 _640_ (.A(net113),
    .B(_307_),
    .Y(_311_));
 sky130_fd_sc_hd__xor2_1 _641_ (.A(\dll_control.tval[1] ),
    .B(_307_),
    .X(_312_));
 sky130_fd_sc_hd__and2_1 _642_ (.A(\dll_control.tval[1] ),
    .B(_307_),
    .X(_313_));
 sky130_fd_sc_hd__a21oi_1 _643_ (.A1(\dll_control.tval[0] ),
    .A2(_312_),
    .B1(_313_),
    .Y(_314_));
 sky130_fd_sc_hd__xnor2_1 _644_ (.A(\dll_control.tval[2] ),
    .B(_307_),
    .Y(_315_));
 sky130_fd_sc_hd__nand2_1 _645_ (.A(\dll_control.tval[2] ),
    .B(_307_),
    .Y(_316_));
 sky130_fd_sc_hd__o21a_1 _646_ (.A1(_314_),
    .A2(_315_),
    .B1(_316_),
    .X(_317_));
 sky130_fd_sc_hd__and2_1 _647_ (.A(net113),
    .B(_307_),
    .X(_318_));
 sky130_fd_sc_hd__o21ba_1 _648_ (.A1(_311_),
    .A2(_317_),
    .B1_N(_318_),
    .X(_319_));
 sky130_fd_sc_hd__and2_1 _649_ (.A(net111),
    .B(_308_),
    .X(_320_));
 sky130_fd_sc_hd__o21ba_1 _650_ (.A1(_310_),
    .A2(_319_),
    .B1_N(_320_),
    .X(_321_));
 sky130_fd_sc_hd__nand2_1 _651_ (.A(net110),
    .B(_308_),
    .Y(_322_));
 sky130_fd_sc_hd__o21ai_1 _652_ (.A1(_309_),
    .A2(_321_),
    .B1(_322_),
    .Y(_323_));
 sky130_fd_sc_hd__nand2b_1 _653_ (.A_N(\dll_control.accum[0] ),
    .B(div[0]),
    .Y(_324_));
 sky130_fd_sc_hd__and4b_1 _654_ (.A_N(_303_),
    .B(_301_),
    .C(_302_),
    .D(_324_),
    .X(_325_));
 sky130_fd_sc_hd__a31o_1 _655_ (.A1(_295_),
    .A2(_300_),
    .A3(_325_),
    .B1(_216_),
    .X(_326_));
 sky130_fd_sc_hd__and3_1 _656_ (.A(\dll_control.tval[2] ),
    .B(\dll_control.tval[1] ),
    .C(\dll_control.tval[0] ),
    .X(_327_));
 sky130_fd_sc_hd__and2_1 _657_ (.A(net112),
    .B(net113),
    .X(_328_));
 sky130_fd_sc_hd__a41o_1 _658_ (.A1(net108),
    .A2(net110),
    .A3(_327_),
    .A4(_328_),
    .B1(net107),
    .X(_329_));
 sky130_fd_sc_hd__nand2b_1 _659_ (.A_N(_308_),
    .B(_329_),
    .Y(_330_));
 sky130_fd_sc_hd__nor2_1 _660_ (.A(net109),
    .B(\dll_control.tint[2] ),
    .Y(_331_));
 sky130_fd_sc_hd__nor2b_1 _661_ (.A(net104),
    .B_N(_331_),
    .Y(_332_));
 sky130_fd_sc_hd__nor2_2 _662_ (.A(net111),
    .B(net113),
    .Y(_333_));
 sky130_fd_sc_hd__nand2_1 _663_ (.A(_332_),
    .B(_333_),
    .Y(_334_));
 sky130_fd_sc_hd__nor3_1 _664_ (.A(\dll_control.tval[1] ),
    .B(\dll_control.tval[0] ),
    .C(_334_),
    .Y(_335_));
 sky130_fd_sc_hd__nand3b_1 _665_ (.A_N(\dll_control.tval[2] ),
    .B(_308_),
    .C(_335_),
    .Y(_336_));
 sky130_fd_sc_hd__nand3b_2 _666_ (.A_N(_326_),
    .B(_330_),
    .C(_336_),
    .Y(_337_));
 sky130_fd_sc_hd__clkbuf_2 _667_ (.A(_337_),
    .X(_338_));
 sky130_fd_sc_hd__o31a_1 _668_ (.A1(net108),
    .A2(_323_),
    .A3(_338_),
    .B1(net106),
    .X(_081_));
 sky130_fd_sc_hd__xnor2_1 _669_ (.A(net108),
    .B(_308_),
    .Y(_339_));
 sky130_fd_sc_hd__xnor2_1 _670_ (.A(_323_),
    .B(_339_),
    .Y(_340_));
 sky130_fd_sc_hd__mux2_1 _671_ (.A0(_340_),
    .A1(net108),
    .S(_338_),
    .X(_341_));
 sky130_fd_sc_hd__clkbuf_1 _672_ (.A(_341_),
    .X(_080_));
 sky130_fd_sc_hd__and2b_1 _673_ (.A_N(_309_),
    .B(_322_),
    .X(_342_));
 sky130_fd_sc_hd__xnor2_1 _674_ (.A(_321_),
    .B(_342_),
    .Y(_343_));
 sky130_fd_sc_hd__mux2_1 _675_ (.A0(_343_),
    .A1(net110),
    .S(_337_),
    .X(_344_));
 sky130_fd_sc_hd__clkbuf_1 _676_ (.A(_344_),
    .X(_079_));
 sky130_fd_sc_hd__nor2_1 _677_ (.A(_320_),
    .B(_310_),
    .Y(_345_));
 sky130_fd_sc_hd__xnor2_1 _678_ (.A(_345_),
    .B(_319_),
    .Y(_346_));
 sky130_fd_sc_hd__mux2_1 _679_ (.A0(_346_),
    .A1(net111),
    .S(_337_),
    .X(_347_));
 sky130_fd_sc_hd__clkbuf_1 _680_ (.A(_347_),
    .X(_078_));
 sky130_fd_sc_hd__nor2_1 _681_ (.A(_311_),
    .B(_318_),
    .Y(_348_));
 sky130_fd_sc_hd__xnor2_1 _682_ (.A(_317_),
    .B(_348_),
    .Y(_349_));
 sky130_fd_sc_hd__mux2_1 _683_ (.A0(_349_),
    .A1(net113),
    .S(_337_),
    .X(_350_));
 sky130_fd_sc_hd__clkbuf_1 _684_ (.A(_350_),
    .X(_077_));
 sky130_fd_sc_hd__xnor2_1 _685_ (.A(_314_),
    .B(_315_),
    .Y(_351_));
 sky130_fd_sc_hd__nor2_1 _686_ (.A(_338_),
    .B(_351_),
    .Y(_352_));
 sky130_fd_sc_hd__a21o_1 _687_ (.A1(\dll_control.tval[2] ),
    .A2(_338_),
    .B1(_352_),
    .X(_076_));
 sky130_fd_sc_hd__nor2_1 _688_ (.A(\dll_control.tval[0] ),
    .B(_312_),
    .Y(_353_));
 sky130_fd_sc_hd__a211o_1 _689_ (.A1(\dll_control.tval[0] ),
    .A2(_312_),
    .B1(_338_),
    .C1(_353_),
    .X(_354_));
 sky130_fd_sc_hd__a21bo_1 _690_ (.A1(\dll_control.tval[1] ),
    .A2(_338_),
    .B1_N(_354_),
    .X(_075_));
 sky130_fd_sc_hd__xnor2_1 _691_ (.A(\dll_control.tval[0] ),
    .B(_338_),
    .Y(_074_));
 sky130_fd_sc_hd__mux2_1 _692_ (.A0(_334_),
    .A1(ext_trim[0]),
    .S(net119),
    .X(_355_));
 sky130_fd_sc_hd__clkbuf_1 _693_ (.A(_355_),
    .X(\itrim[0] ));
 sky130_fd_sc_hd__inv_2 _694_ (.A(_333_),
    .Y(_356_));
 sky130_fd_sc_hd__nand2_1 _695_ (.A(net112),
    .B(net113),
    .Y(_357_));
 sky130_fd_sc_hd__and2b_1 _696_ (.A_N(net109),
    .B(net110),
    .X(_358_));
 sky130_fd_sc_hd__and2b_1 _697_ (.A_N(net104),
    .B(_358_),
    .X(_359_));
 sky130_fd_sc_hd__nand3_1 _698_ (.A(_356_),
    .B(_357_),
    .C(_359_),
    .Y(_360_));
 sky130_fd_sc_hd__nand2_1 _699_ (.A(_333_),
    .B(_359_),
    .Y(_361_));
 sky130_fd_sc_hd__nor2_2 _700_ (.A(net122),
    .B(_332_),
    .Y(_362_));
 sky130_fd_sc_hd__and3_1 _701_ (.A(_360_),
    .B(_361_),
    .C(_362_),
    .X(_363_));
 sky130_fd_sc_hd__and2b_1 _702_ (.A_N(net110),
    .B(net108),
    .X(_364_));
 sky130_fd_sc_hd__a22o_1 _703_ (.A1(_328_),
    .A2(_358_),
    .B1(_364_),
    .B2(_333_),
    .X(_365_));
 sky130_fd_sc_hd__nand2b_1 _704_ (.A_N(net105),
    .B(_365_),
    .Y(_366_));
 sky130_fd_sc_hd__nand3b_1 _705_ (.A_N(net104),
    .B(_356_),
    .C(_364_),
    .Y(_367_));
 sky130_fd_sc_hd__and3_1 _706_ (.A(_363_),
    .B(_366_),
    .C(_367_),
    .X(_368_));
 sky130_fd_sc_hd__a21o_1 _707_ (.A1(net119),
    .A2(ext_trim[1]),
    .B1(_368_),
    .X(\itrim[1] ));
 sky130_fd_sc_hd__o21ba_1 _708_ (.A1(net107),
    .A2(net108),
    .B1_N(net122),
    .X(_369_));
 sky130_fd_sc_hd__a21o_1 _709_ (.A1(net119),
    .A2(ext_trim[2]),
    .B1(_369_),
    .X(\itrim[2] ));
 sky130_fd_sc_hd__a21o_1 _710_ (.A1(net118),
    .A2(ext_trim[3]),
    .B1(_362_),
    .X(\itrim[3] ));
 sky130_fd_sc_hd__nand2_1 _711_ (.A(\dll_control.tint[0] ),
    .B(_364_),
    .Y(_370_));
 sky130_fd_sc_hd__and2_1 _712_ (.A(_363_),
    .B(_366_),
    .X(_371_));
 sky130_fd_sc_hd__o31a_1 _713_ (.A1(net107),
    .A2(net111),
    .A3(_370_),
    .B1(_371_),
    .X(_372_));
 sky130_fd_sc_hd__a21o_1 _714_ (.A1(net118),
    .A2(ext_trim[4]),
    .B1(_372_),
    .X(\itrim[4] ));
 sky130_fd_sc_hd__a21o_1 _715_ (.A1(net118),
    .A2(ext_trim[5]),
    .B1(_363_),
    .X(\itrim[5] ));
 sky130_fd_sc_hd__mux2_1 _716_ (.A0(net111),
    .A1(ext_trim[6]),
    .S(net118),
    .X(_373_));
 sky130_fd_sc_hd__nor2_1 _717_ (.A(_362_),
    .B(_373_),
    .Y(_374_));
 sky130_fd_sc_hd__inv_2 _718_ (.A(_374_),
    .Y(\itrim[6] ));
 sky130_fd_sc_hd__nand3b_2 _719_ (.A_N(net104),
    .B(net108),
    .C(net110),
    .Y(_375_));
 sky130_fd_sc_hd__and2_1 _720_ (.A(_368_),
    .B(_375_),
    .X(_376_));
 sky130_fd_sc_hd__clkbuf_2 _721_ (.A(_376_),
    .X(_377_));
 sky130_fd_sc_hd__a221o_1 _722_ (.A1(net121),
    .A2(ext_trim[7]),
    .B1(_356_),
    .B2(_368_),
    .C1(_377_),
    .X(\itrim[7] ));
 sky130_fd_sc_hd__a22o_1 _723_ (.A1(net120),
    .A2(ext_trim[8]),
    .B1(_361_),
    .B2(_362_),
    .X(\itrim[8] ));
 sky130_fd_sc_hd__a21o_1 _724_ (.A1(net122),
    .A2(ext_trim[9]),
    .B1(_371_),
    .X(\itrim[9] ));
 sky130_fd_sc_hd__a21oi_1 _725_ (.A1(_332_),
    .A2(_357_),
    .B1(net120),
    .Y(_378_));
 sky130_fd_sc_hd__a21o_1 _726_ (.A1(net121),
    .A2(ext_trim[10]),
    .B1(_378_),
    .X(\itrim[10] ));
 sky130_fd_sc_hd__a221o_2 _727_ (.A1(net120),
    .A2(ext_trim[11]),
    .B1(_328_),
    .B2(_371_),
    .C1(_368_),
    .X(\itrim[11] ));
 sky130_fd_sc_hd__inv_2 _728_ (.A(net112),
    .Y(_379_));
 sky130_fd_sc_hd__nand2_1 _729_ (.A(_379_),
    .B(_359_),
    .Y(_380_));
 sky130_fd_sc_hd__a22o_1 _730_ (.A1(net120),
    .A2(ext_trim[12]),
    .B1(_380_),
    .B2(_362_),
    .X(\itrim[12] ));
 sky130_fd_sc_hd__o21a_1 _731_ (.A1(net111),
    .A2(_375_),
    .B1(_368_),
    .X(_381_));
 sky130_fd_sc_hd__a21o_1 _732_ (.A1(net120),
    .A2(ext_trim[13]),
    .B1(_381_),
    .X(\itrim[13] ));
 sky130_fd_sc_hd__nand2_1 _733_ (.A(_332_),
    .B(_328_),
    .Y(_382_));
 sky130_fd_sc_hd__and4_1 _734_ (.A(_360_),
    .B(_361_),
    .C(_382_),
    .D(_367_),
    .X(_383_));
 sky130_fd_sc_hd__and3b_1 _735_ (.A_N(net120),
    .B(_375_),
    .C(_383_),
    .X(_384_));
 sky130_fd_sc_hd__and2_1 _736_ (.A(net105),
    .B(_358_),
    .X(_385_));
 sky130_fd_sc_hd__nand2_1 _737_ (.A(_357_),
    .B(_385_),
    .Y(_386_));
 sky130_fd_sc_hd__nand2_1 _738_ (.A(net105),
    .B(_331_),
    .Y(_387_));
 sky130_fd_sc_hd__nand2_1 _739_ (.A(_331_),
    .B(_357_),
    .Y(_388_));
 sky130_fd_sc_hd__and4b_1 _740_ (.A_N(_365_),
    .B(_386_),
    .C(_387_),
    .D(_388_),
    .X(_389_));
 sky130_fd_sc_hd__a22o_1 _741_ (.A1(net135),
    .A2(ext_trim[14]),
    .B1(_384_),
    .B2(_389_),
    .X(\itrim[14] ));
 sky130_fd_sc_hd__and3_1 _742_ (.A(_368_),
    .B(_375_),
    .C(_387_),
    .X(_390_));
 sky130_fd_sc_hd__nand2_1 _743_ (.A(_333_),
    .B(_385_),
    .Y(_391_));
 sky130_fd_sc_hd__a22o_1 _744_ (.A1(net135),
    .A2(ext_trim[15]),
    .B1(_390_),
    .B2(_391_),
    .X(\itrim[15] ));
 sky130_fd_sc_hd__nand2_1 _745_ (.A(_331_),
    .B(_333_),
    .Y(_392_));
 sky130_fd_sc_hd__a22o_1 _746_ (.A1(net135),
    .A2(ext_trim[16]),
    .B1(_377_),
    .B2(_392_),
    .X(\itrim[16] ));
 sky130_fd_sc_hd__a22o_1 _747_ (.A1(net135),
    .A2(ext_trim[17]),
    .B1(_386_),
    .B2(_390_),
    .X(\itrim[17] ));
 sky130_fd_sc_hd__a21o_1 _748_ (.A1(net136),
    .A2(ext_trim[18]),
    .B1(_390_),
    .X(\itrim[18] ));
 sky130_fd_sc_hd__o211a_1 _749_ (.A1(_328_),
    .A2(_375_),
    .B1(_366_),
    .C1(_378_),
    .X(_393_));
 sky130_fd_sc_hd__a22o_1 _750_ (.A1(net120),
    .A2(ext_trim[19]),
    .B1(_383_),
    .B2(_393_),
    .X(\itrim[19] ));
 sky130_fd_sc_hd__nand4_1 _751_ (.A(net105),
    .B(_379_),
    .C(net113),
    .D(_364_),
    .Y(_394_));
 sky130_fd_sc_hd__a32o_1 _752_ (.A1(_384_),
    .A2(_389_),
    .A3(_394_),
    .B1(ext_trim[20]),
    .B2(net135),
    .X(\itrim[20] ));
 sky130_fd_sc_hd__nand2b_1 _753_ (.A_N(net104),
    .B(_331_),
    .Y(_395_));
 sky130_fd_sc_hd__o22a_1 _754_ (.A1(_395_),
    .A2(_328_),
    .B1(_387_),
    .B2(net112),
    .X(_396_));
 sky130_fd_sc_hd__a32o_1 _755_ (.A1(_366_),
    .A2(_384_),
    .A3(_396_),
    .B1(ext_trim[21]),
    .B2(net135),
    .X(\itrim[21] ));
 sky130_fd_sc_hd__a31o_1 _756_ (.A1(net104),
    .A2(_379_),
    .A3(_358_),
    .B1(_331_),
    .X(_397_));
 sky130_fd_sc_hd__o21ai_1 _757_ (.A1(net104),
    .A2(_357_),
    .B1(_397_),
    .Y(_398_));
 sky130_fd_sc_hd__a32o_1 _758_ (.A1(_366_),
    .A2(_384_),
    .A3(_398_),
    .B1(ext_trim[22]),
    .B2(net135),
    .X(\itrim[22] ));
 sky130_fd_sc_hd__a21o_1 _759_ (.A1(net137),
    .A2(ext_trim[23]),
    .B1(_377_),
    .X(\itrim[23] ));
 sky130_fd_sc_hd__a22o_1 _760_ (.A1(net137),
    .A2(ext_trim[24]),
    .B1(_377_),
    .B2(net109),
    .X(\itrim[24] ));
 sky130_fd_sc_hd__a22o_1 _761_ (.A1(net136),
    .A2(ext_trim[25]),
    .B1(_388_),
    .B2(_377_),
    .X(\itrim[25] ));
 sky130_fd_sc_hd__nand2_1 _762_ (.A(enable),
    .B(resetb),
    .Y(_399_));
 sky130_fd_sc_hd__clkbuf_1 _763_ (.A(_399_),
    .X(ireset));
 sky130_fd_sc_hd__nor2_1 _764_ (.A(net118),
    .B(net114),
    .Y(_000_));
 sky130_fd_sc_hd__nor2_1 _765_ (.A(net118),
    .B(net114),
    .Y(_001_));
 sky130_fd_sc_hd__nor2_1 _766_ (.A(net118),
    .B(net114),
    .Y(_002_));
 sky130_fd_sc_hd__nor2_1 _767_ (.A(net123),
    .B(ireset),
    .Y(_003_));
 sky130_fd_sc_hd__nor2_1 _768_ (.A(net123),
    .B(net114),
    .Y(_004_));
 sky130_fd_sc_hd__nor2_1 _769_ (.A(net123),
    .B(net114),
    .Y(_005_));
 sky130_fd_sc_hd__clkbuf_2 _770_ (.A(_399_),
    .X(_400_));
 sky130_fd_sc_hd__clkbuf_2 _771_ (.A(_400_),
    .X(_401_));
 sky130_fd_sc_hd__nor2_1 _772_ (.A(net137),
    .B(_401_),
    .Y(_006_));
 sky130_fd_sc_hd__nor2_1 _773_ (.A(net137),
    .B(_401_),
    .Y(_007_));
 sky130_fd_sc_hd__nor2_1 _774_ (.A(net137),
    .B(_401_),
    .Y(_008_));
 sky130_fd_sc_hd__nor2_1 _775_ (.A(net137),
    .B(_401_),
    .Y(_009_));
 sky130_fd_sc_hd__nor2_1 _776_ (.A(net137),
    .B(_401_),
    .Y(_010_));
 sky130_fd_sc_hd__nor2_1 _777_ (.A(net138),
    .B(_401_),
    .Y(_011_));
 sky130_fd_sc_hd__nor2_1 _778_ (.A(net138),
    .B(_401_),
    .Y(_012_));
 sky130_fd_sc_hd__clkbuf_2 _779_ (.A(_400_),
    .X(_402_));
 sky130_fd_sc_hd__nor2_1 _780_ (.A(net132),
    .B(_402_),
    .Y(_013_));
 sky130_fd_sc_hd__nor2_1 _781_ (.A(net129),
    .B(_402_),
    .Y(_014_));
 sky130_fd_sc_hd__nor2_1 _782_ (.A(net130),
    .B(_402_),
    .Y(_015_));
 sky130_fd_sc_hd__nor2_1 _783_ (.A(net130),
    .B(_402_),
    .Y(_016_));
 sky130_fd_sc_hd__nor2_1 _784_ (.A(net130),
    .B(_402_),
    .Y(_017_));
 sky130_fd_sc_hd__nor2_1 _785_ (.A(net130),
    .B(_402_),
    .Y(_018_));
 sky130_fd_sc_hd__nor2_1 _786_ (.A(net132),
    .B(_402_),
    .Y(_019_));
 sky130_fd_sc_hd__clkbuf_2 _787_ (.A(_399_),
    .X(_403_));
 sky130_fd_sc_hd__clkbuf_2 _788_ (.A(_403_),
    .X(_404_));
 sky130_fd_sc_hd__nor2_1 _789_ (.A(net116),
    .B(_404_),
    .Y(_020_));
 sky130_fd_sc_hd__nor2_1 _790_ (.A(net127),
    .B(_404_),
    .Y(_021_));
 sky130_fd_sc_hd__nor2_1 _791_ (.A(net127),
    .B(_404_),
    .Y(_022_));
 sky130_fd_sc_hd__nor2_1 _792_ (.A(net127),
    .B(_404_),
    .Y(_023_));
 sky130_fd_sc_hd__nor2_1 _793_ (.A(net127),
    .B(_404_),
    .Y(_024_));
 sky130_fd_sc_hd__nor2_1 _794_ (.A(net128),
    .B(_404_),
    .Y(_025_));
 sky130_fd_sc_hd__nor2_1 _795_ (.A(net127),
    .B(_404_),
    .Y(_026_));
 sky130_fd_sc_hd__clkbuf_2 _796_ (.A(_403_),
    .X(_405_));
 sky130_fd_sc_hd__nor2_1 _797_ (.A(net131),
    .B(_405_),
    .Y(_027_));
 sky130_fd_sc_hd__nor2_1 _798_ (.A(net131),
    .B(_405_),
    .Y(_028_));
 sky130_fd_sc_hd__nor2_1 _799_ (.A(net130),
    .B(_405_),
    .Y(_029_));
 sky130_fd_sc_hd__nor2_1 _800_ (.A(net131),
    .B(_405_),
    .Y(_030_));
 sky130_fd_sc_hd__nor2_1 _801_ (.A(net131),
    .B(_405_),
    .Y(_031_));
 sky130_fd_sc_hd__nor2_1 _802_ (.A(net116),
    .B(_405_),
    .Y(_032_));
 sky130_fd_sc_hd__nor2_1 _803_ (.A(net116),
    .B(_405_),
    .Y(_033_));
 sky130_fd_sc_hd__clkbuf_2 _804_ (.A(_403_),
    .X(_406_));
 sky130_fd_sc_hd__nor2_1 _805_ (.A(net117),
    .B(_406_),
    .Y(_034_));
 sky130_fd_sc_hd__nor2_1 _806_ (.A(net117),
    .B(_406_),
    .Y(_035_));
 sky130_fd_sc_hd__nor2_1 _807_ (.A(net116),
    .B(_406_),
    .Y(_036_));
 sky130_fd_sc_hd__nor2_1 _808_ (.A(net117),
    .B(_406_),
    .Y(_037_));
 sky130_fd_sc_hd__nor2_1 _809_ (.A(net126),
    .B(_406_),
    .Y(_038_));
 sky130_fd_sc_hd__nor2_1 _810_ (.A(net126),
    .B(_406_),
    .Y(_039_));
 sky130_fd_sc_hd__nor2_1 _811_ (.A(net126),
    .B(_406_),
    .Y(_040_));
 sky130_fd_sc_hd__clkbuf_2 _812_ (.A(_403_),
    .X(_407_));
 sky130_fd_sc_hd__nor2_1 _813_ (.A(net128),
    .B(_407_),
    .Y(_041_));
 sky130_fd_sc_hd__nor2_1 _814_ (.A(net132),
    .B(_407_),
    .Y(_042_));
 sky130_fd_sc_hd__nor2_1 _815_ (.A(net133),
    .B(_407_),
    .Y(_043_));
 sky130_fd_sc_hd__nor2_1 _816_ (.A(net128),
    .B(_407_),
    .Y(_044_));
 sky130_fd_sc_hd__nor2_1 _817_ (.A(net132),
    .B(_407_),
    .Y(_045_));
 sky130_fd_sc_hd__nor2_1 _818_ (.A(net132),
    .B(_407_),
    .Y(_046_));
 sky130_fd_sc_hd__nor2_1 _819_ (.A(net133),
    .B(_407_),
    .Y(_047_));
 sky130_fd_sc_hd__buf_2 _820_ (.A(_403_),
    .X(_408_));
 sky130_fd_sc_hd__nor2_1 _821_ (.A(net133),
    .B(_408_),
    .Y(_048_));
 sky130_fd_sc_hd__nor2_1 _822_ (.A(net133),
    .B(_408_),
    .Y(_049_));
 sky130_fd_sc_hd__nor2_1 _823_ (.A(net130),
    .B(_408_),
    .Y(_050_));
 sky130_fd_sc_hd__nor2_1 _824_ (.A(net131),
    .B(_408_),
    .Y(_051_));
 sky130_fd_sc_hd__nor2_1 _825_ (.A(net130),
    .B(_408_),
    .Y(_052_));
 sky130_fd_sc_hd__nor2_1 _826_ (.A(net126),
    .B(_408_),
    .Y(_053_));
 sky130_fd_sc_hd__nor2_1 _827_ (.A(net126),
    .B(_408_),
    .Y(_054_));
 sky130_fd_sc_hd__clkbuf_2 _828_ (.A(_403_),
    .X(_409_));
 sky130_fd_sc_hd__nor2_1 _829_ (.A(net126),
    .B(_409_),
    .Y(_055_));
 sky130_fd_sc_hd__nor2_1 _830_ (.A(net126),
    .B(_409_),
    .Y(_056_));
 sky130_fd_sc_hd__nor2_1 _831_ (.A(net127),
    .B(_409_),
    .Y(_057_));
 sky130_fd_sc_hd__nor2_1 _832_ (.A(net127),
    .B(_409_),
    .Y(_058_));
 sky130_fd_sc_hd__nor2_1 _833_ (.A(net128),
    .B(_409_),
    .Y(_059_));
 sky130_fd_sc_hd__nor2_1 _834_ (.A(net132),
    .B(_409_),
    .Y(_060_));
 sky130_fd_sc_hd__nor2_1 _835_ (.A(net132),
    .B(_409_),
    .Y(_061_));
 sky130_fd_sc_hd__buf_2 _836_ (.A(_403_),
    .X(_410_));
 sky130_fd_sc_hd__nor2_1 _837_ (.A(net133),
    .B(_410_),
    .Y(_062_));
 sky130_fd_sc_hd__nor2_1 _838_ (.A(net131),
    .B(_410_),
    .Y(_063_));
 sky130_fd_sc_hd__nor2_1 _839_ (.A(net133),
    .B(_410_),
    .Y(_064_));
 sky130_fd_sc_hd__nor2_1 _840_ (.A(net115),
    .B(_410_),
    .Y(_065_));
 sky130_fd_sc_hd__nor2_1 _841_ (.A(net115),
    .B(_410_),
    .Y(_066_));
 sky130_fd_sc_hd__nor2_1 _842_ (.A(net115),
    .B(_410_),
    .Y(_067_));
 sky130_fd_sc_hd__nor2_1 _843_ (.A(net115),
    .B(_410_),
    .Y(_068_));
 sky130_fd_sc_hd__nor2_1 _844_ (.A(net116),
    .B(_400_),
    .Y(_069_));
 sky130_fd_sc_hd__nor2_1 _845_ (.A(net116),
    .B(_400_),
    .Y(_070_));
 sky130_fd_sc_hd__nor2_1 _846_ (.A(net115),
    .B(_400_),
    .Y(_071_));
 sky130_fd_sc_hd__nor2_1 _847_ (.A(net115),
    .B(_400_),
    .Y(_072_));
 sky130_fd_sc_hd__nor2_1 _848_ (.A(net115),
    .B(_400_),
    .Y(_073_));
 sky130_fd_sc_hd__dfrtp_1 _849_ (.CLK(\clockp_buffer_in[0] ),
    .D(_074_),
    .RESET_B(_000_),
    .Q(\dll_control.tval[0] ));
 sky130_fd_sc_hd__dfrtp_1 _850_ (.CLK(\clockp_buffer_in[0] ),
    .D(_075_),
    .RESET_B(_001_),
    .Q(\dll_control.tval[1] ));
 sky130_fd_sc_hd__dfrtp_1 _851_ (.CLK(\clockp_buffer_in[0] ),
    .D(_076_),
    .RESET_B(_002_),
    .Q(\dll_control.tval[2] ));
 sky130_fd_sc_hd__dfrtp_1 _852_ (.CLK(\clockp_buffer_in[0] ),
    .D(_077_),
    .RESET_B(_003_),
    .Q(\dll_control.tint[0] ));
 sky130_fd_sc_hd__dfrtp_1 _853_ (.CLK(\clockp_buffer_in[0] ),
    .D(_078_),
    .RESET_B(_004_),
    .Q(\dll_control.tint[1] ));
 sky130_fd_sc_hd__dfrtp_1 _854_ (.CLK(\clockp_buffer_in[0] ),
    .D(_079_),
    .RESET_B(_005_),
    .Q(\dll_control.tint[2] ));
 sky130_fd_sc_hd__dfrtp_1 _855_ (.CLK(\clockp_buffer_in[0] ),
    .D(_080_),
    .RESET_B(_006_),
    .Q(\dll_control.tint[3] ));
 sky130_fd_sc_hd__dfrtp_1 _856_ (.CLK(\clockp_buffer_in[0] ),
    .D(_081_),
    .RESET_B(_007_),
    .Q(\dll_control.tint[4] ));
 sky130_fd_sc_hd__dfrtp_1 _857_ (.CLK(\clockp_buffer_in[0] ),
    .D(_082_),
    .RESET_B(_008_),
    .Q(\dll_control.count2[0] ));
 sky130_fd_sc_hd__dfrtp_1 _858_ (.CLK(\clockp_buffer_in[0] ),
    .D(_083_),
    .RESET_B(_009_),
    .Q(\dll_control.count2[1] ));
 sky130_fd_sc_hd__dfrtp_1 _859_ (.CLK(\clockp_buffer_in[0] ),
    .D(_084_),
    .RESET_B(_010_),
    .Q(\dll_control.count2[2] ));
 sky130_fd_sc_hd__dfrtp_1 _860_ (.CLK(\clockp_buffer_in[0] ),
    .D(_085_),
    .RESET_B(_011_),
    .Q(\dll_control.count2[3] ));
 sky130_fd_sc_hd__dfrtp_1 _861_ (.CLK(\clockp_buffer_in[0] ),
    .D(_086_),
    .RESET_B(_012_),
    .Q(\dll_control.count2[4] ));
 sky130_fd_sc_hd__dfrtp_1 _862_ (.CLK(\clockp_buffer_in[0] ),
    .D(_087_),
    .RESET_B(_013_),
    .Q(\dll_control.count2[5] ));
 sky130_fd_sc_hd__dfrtp_1 _863_ (.CLK(\clockp_buffer_in[0] ),
    .D(_088_),
    .RESET_B(_014_),
    .Q(\dll_control.count6[0] ));
 sky130_fd_sc_hd__dfrtp_1 _864_ (.CLK(\clockp_buffer_in[0] ),
    .D(_089_),
    .RESET_B(_015_),
    .Q(\dll_control.count6[1] ));
 sky130_fd_sc_hd__dfrtp_1 _865_ (.CLK(\clockp_buffer_in[0] ),
    .D(_090_),
    .RESET_B(_016_),
    .Q(\dll_control.count6[2] ));
 sky130_fd_sc_hd__dfrtp_1 _866_ (.CLK(\clockp_buffer_in[0] ),
    .D(_091_),
    .RESET_B(_017_),
    .Q(\dll_control.count6[3] ));
 sky130_fd_sc_hd__dfrtp_1 _867_ (.CLK(\clockp_buffer_in[0] ),
    .D(_092_),
    .RESET_B(_018_),
    .Q(\dll_control.count6[4] ));
 sky130_fd_sc_hd__dfrtp_1 _868_ (.CLK(\clockp_buffer_in[0] ),
    .D(_093_),
    .RESET_B(_019_),
    .Q(\dll_control.count6[5] ));
 sky130_fd_sc_hd__dfrtp_1 _869_ (.CLK(\clockp_buffer_in[0] ),
    .D(_094_),
    .RESET_B(_020_),
    .Q(\dll_control.count1[0] ));
 sky130_fd_sc_hd__dfrtp_1 _870_ (.CLK(\clockp_buffer_in[0] ),
    .D(_095_),
    .RESET_B(_021_),
    .Q(\dll_control.count1[1] ));
 sky130_fd_sc_hd__dfrtp_1 _871_ (.CLK(\clockp_buffer_in[0] ),
    .D(_096_),
    .RESET_B(_022_),
    .Q(\dll_control.count1[2] ));
 sky130_fd_sc_hd__dfrtp_1 _872_ (.CLK(\clockp_buffer_in[0] ),
    .D(_097_),
    .RESET_B(_023_),
    .Q(\dll_control.count1[3] ));
 sky130_fd_sc_hd__dfrtp_1 _873_ (.CLK(\clockp_buffer_in[0] ),
    .D(_098_),
    .RESET_B(_024_),
    .Q(\dll_control.count1[4] ));
 sky130_fd_sc_hd__dfrtp_1 _874_ (.CLK(\clockp_buffer_in[0] ),
    .D(_099_),
    .RESET_B(_025_),
    .Q(\dll_control.count1[5] ));
 sky130_fd_sc_hd__dfrtp_1 _875_ (.CLK(\clockp_buffer_in[0] ),
    .D(_100_),
    .RESET_B(_026_),
    .Q(\dll_control.count5[0] ));
 sky130_fd_sc_hd__dfrtp_1 _876_ (.CLK(\clockp_buffer_in[0] ),
    .D(_101_),
    .RESET_B(_027_),
    .Q(\dll_control.count5[1] ));
 sky130_fd_sc_hd__dfrtp_1 _877_ (.CLK(\clockp_buffer_in[0] ),
    .D(_102_),
    .RESET_B(_028_),
    .Q(\dll_control.count5[2] ));
 sky130_fd_sc_hd__dfrtp_1 _878_ (.CLK(\clockp_buffer_in[0] ),
    .D(_103_),
    .RESET_B(_029_),
    .Q(\dll_control.count5[3] ));
 sky130_fd_sc_hd__dfrtp_1 _879_ (.CLK(\clockp_buffer_in[0] ),
    .D(_104_),
    .RESET_B(_030_),
    .Q(\dll_control.count5[4] ));
 sky130_fd_sc_hd__dfrtp_1 _880_ (.CLK(\clockp_buffer_in[0] ),
    .D(_105_),
    .RESET_B(_031_),
    .Q(\dll_control.count5[5] ));
 sky130_fd_sc_hd__dfrtp_2 _881_ (.CLK(\clockp_buffer_in[0] ),
    .D(_106_),
    .RESET_B(_032_),
    .Q(\dll_control.count0[0] ));
 sky130_fd_sc_hd__dfrtp_2 _882_ (.CLK(\clockp_buffer_in[0] ),
    .D(_107_),
    .RESET_B(_033_),
    .Q(\dll_control.count0[1] ));
 sky130_fd_sc_hd__dfrtp_1 _883_ (.CLK(\clockp_buffer_in[0] ),
    .D(_108_),
    .RESET_B(_034_),
    .Q(\dll_control.count0[2] ));
 sky130_fd_sc_hd__dfrtp_2 _884_ (.CLK(\clockp_buffer_in[0] ),
    .D(_109_),
    .RESET_B(_035_),
    .Q(\dll_control.count0[3] ));
 sky130_fd_sc_hd__dfrtp_1 _885_ (.CLK(\clockp_buffer_in[0] ),
    .D(_110_),
    .RESET_B(_036_),
    .Q(\dll_control.count0[4] ));
 sky130_fd_sc_hd__dfrtp_1 _886_ (.CLK(\clockp_buffer_in[0] ),
    .D(_111_),
    .RESET_B(_037_),
    .Q(\dll_control.count0[5] ));
 sky130_fd_sc_hd__dfrtp_1 _887_ (.CLK(\clockp_buffer_in[0] ),
    .D(_112_),
    .RESET_B(_038_),
    .Q(\dll_control.count7[0] ));
 sky130_fd_sc_hd__dfrtp_1 _888_ (.CLK(\clockp_buffer_in[0] ),
    .D(_113_),
    .RESET_B(_039_),
    .Q(\dll_control.count7[1] ));
 sky130_fd_sc_hd__dfrtp_1 _889_ (.CLK(\clockp_buffer_in[0] ),
    .D(_114_),
    .RESET_B(_040_),
    .Q(\dll_control.count7[2] ));
 sky130_fd_sc_hd__dfrtp_1 _890_ (.CLK(\clockp_buffer_in[0] ),
    .D(_115_),
    .RESET_B(_041_),
    .Q(\dll_control.count7[3] ));
 sky130_fd_sc_hd__dfrtp_1 _891_ (.CLK(\clockp_buffer_in[0] ),
    .D(_116_),
    .RESET_B(_042_),
    .Q(\dll_control.count7[4] ));
 sky130_fd_sc_hd__dfrtp_1 _892_ (.CLK(\clockp_buffer_in[0] ),
    .D(_117_),
    .RESET_B(_043_),
    .Q(\dll_control.count7[5] ));
 sky130_fd_sc_hd__dfrtp_1 _893_ (.CLK(\clockp_buffer_in[0] ),
    .D(_118_),
    .RESET_B(_044_),
    .Q(\dll_control.count3[0] ));
 sky130_fd_sc_hd__dfrtp_1 _894_ (.CLK(\clockp_buffer_in[0] ),
    .D(_119_),
    .RESET_B(_045_),
    .Q(\dll_control.count3[1] ));
 sky130_fd_sc_hd__dfrtp_1 _895_ (.CLK(\clockp_buffer_in[0] ),
    .D(_120_),
    .RESET_B(_046_),
    .Q(\dll_control.count3[2] ));
 sky130_fd_sc_hd__dfrtp_1 _896_ (.CLK(\clockp_buffer_in[0] ),
    .D(_121_),
    .RESET_B(_047_),
    .Q(\dll_control.count3[3] ));
 sky130_fd_sc_hd__dfrtp_1 _897_ (.CLK(\clockp_buffer_in[0] ),
    .D(_122_),
    .RESET_B(_048_),
    .Q(\dll_control.count3[4] ));
 sky130_fd_sc_hd__dfrtp_1 _898_ (.CLK(\clockp_buffer_in[0] ),
    .D(_123_),
    .RESET_B(_049_),
    .Q(\dll_control.count3[5] ));
 sky130_fd_sc_hd__dfrtp_1 _899_ (.CLK(\clockp_buffer_in[0] ),
    .D(osc),
    .RESET_B(_050_),
    .Q(\dll_control.oscbuf[0] ));
 sky130_fd_sc_hd__dfrtp_1 _900_ (.CLK(\clockp_buffer_in[0] ),
    .D(\dll_control.oscbuf[0] ),
    .RESET_B(_051_),
    .Q(\dll_control.oscbuf[1] ));
 sky130_fd_sc_hd__dfrtp_1 _901_ (.CLK(\clockp_buffer_in[0] ),
    .D(\dll_control.oscbuf[1] ),
    .RESET_B(_052_),
    .Q(\dll_control.oscbuf[2] ));
 sky130_fd_sc_hd__dfrtp_1 _902_ (.CLK(\clockp_buffer_in[0] ),
    .D(_124_),
    .RESET_B(_053_),
    .Q(\dll_control.count8[0] ));
 sky130_fd_sc_hd__dfrtp_1 _903_ (.CLK(\clockp_buffer_in[0] ),
    .D(_125_),
    .RESET_B(_054_),
    .Q(\dll_control.count8[1] ));
 sky130_fd_sc_hd__dfrtp_1 _904_ (.CLK(\clockp_buffer_in[0] ),
    .D(_126_),
    .RESET_B(_055_),
    .Q(\dll_control.count8[2] ));
 sky130_fd_sc_hd__dfrtp_1 _905_ (.CLK(\clockp_buffer_in[0] ),
    .D(_127_),
    .RESET_B(_056_),
    .Q(\dll_control.count8[3] ));
 sky130_fd_sc_hd__dfrtp_1 _906_ (.CLK(\clockp_buffer_in[0] ),
    .D(_128_),
    .RESET_B(_057_),
    .Q(\dll_control.count8[4] ));
 sky130_fd_sc_hd__dfrtp_1 _907_ (.CLK(\clockp_buffer_in[0] ),
    .D(_129_),
    .RESET_B(_058_),
    .Q(\dll_control.count8[5] ));
 sky130_fd_sc_hd__dfrtp_1 _908_ (.CLK(\clockp_buffer_in[0] ),
    .D(_130_),
    .RESET_B(_059_),
    .Q(\dll_control.count4[0] ));
 sky130_fd_sc_hd__dfrtp_1 _909_ (.CLK(\clockp_buffer_in[0] ),
    .D(_131_),
    .RESET_B(_060_),
    .Q(\dll_control.count4[1] ));
 sky130_fd_sc_hd__dfrtp_1 _910_ (.CLK(\clockp_buffer_in[0] ),
    .D(_132_),
    .RESET_B(_061_),
    .Q(\dll_control.count4[2] ));
 sky130_fd_sc_hd__dfrtp_1 _911_ (.CLK(\clockp_buffer_in[0] ),
    .D(_133_),
    .RESET_B(_062_),
    .Q(\dll_control.count4[3] ));
 sky130_fd_sc_hd__dfrtp_1 _912_ (.CLK(\clockp_buffer_in[0] ),
    .D(_134_),
    .RESET_B(_063_),
    .Q(\dll_control.count4[4] ));
 sky130_fd_sc_hd__dfrtp_1 _913_ (.CLK(\clockp_buffer_in[0] ),
    .D(_135_),
    .RESET_B(_064_),
    .Q(\dll_control.count4[5] ));
 sky130_fd_sc_hd__dfrtp_1 _914_ (.CLK(\clockp_buffer_in[0] ),
    .D(_136_),
    .RESET_B(_065_),
    .Q(\dll_control.accum[0] ));
 sky130_fd_sc_hd__dfrtp_1 _915_ (.CLK(\clockp_buffer_in[0] ),
    .D(_137_),
    .RESET_B(_066_),
    .Q(\dll_control.accum[1] ));
 sky130_fd_sc_hd__dfrtp_1 _916_ (.CLK(\clockp_buffer_in[0] ),
    .D(_138_),
    .RESET_B(_067_),
    .Q(\dll_control.accum[2] ));
 sky130_fd_sc_hd__dfrtp_1 _917_ (.CLK(\clockp_buffer_in[0] ),
    .D(_139_),
    .RESET_B(_068_),
    .Q(\dll_control.accum[3] ));
 sky130_fd_sc_hd__dfrtp_1 _918_ (.CLK(\clockp_buffer_in[0] ),
    .D(_140_),
    .RESET_B(_069_),
    .Q(\dll_control.accum[4] ));
 sky130_fd_sc_hd__dfrtp_1 _919_ (.CLK(\clockp_buffer_in[0] ),
    .D(_141_),
    .RESET_B(_070_),
    .Q(\dll_control.accum[5] ));
 sky130_fd_sc_hd__dfrtp_1 _920_ (.CLK(\clockp_buffer_in[0] ),
    .D(_142_),
    .RESET_B(_071_),
    .Q(\dll_control.accum[6] ));
 sky130_fd_sc_hd__dfrtp_1 _921_ (.CLK(\clockp_buffer_in[0] ),
    .D(_143_),
    .RESET_B(_072_),
    .Q(\dll_control.accum[7] ));
 sky130_fd_sc_hd__dfrtp_1 _922_ (.CLK(\clockp_buffer_in[0] ),
    .D(_144_),
    .RESET_B(_073_),
    .Q(\dll_control.accum[8] ));
 sky130_fd_sc_hd__clkbuf_16 clockp_buffer_0 (.A(\clockp_buffer_in[0] ),
    .X(clockp[0]));
 sky130_fd_sc_hd__buf_4 clockp_buffer_1 (.A(\clockp_buffer_in[1] ),
    .X(clockp[1]));
 sky130_fd_sc_hd__clkbuf_1 \ringosc.dstage[0].id.delaybuf0  (.A(\ringosc.dstage[0].id.in ),
    .X(\ringosc.dstage[0].id.ts ));
 sky130_fd_sc_hd__clkbuf_1 \ringosc.dstage[0].id.delaybuf1  (.A(\ringosc.dstage[0].id.ts ),
    .X(\ringosc.dstage[0].id.d0 ));
 sky130_fd_sc_hd__einvp_2 \ringosc.dstage[0].id.delayen0  (.A(\ringosc.dstage[0].id.d2 ),
    .TE(\itrim[0] ),
    .Z(\ringosc.dstage[0].id.out ));
 sky130_fd_sc_hd__einvp_1 \ringosc.dstage[0].id.delayen1  (.A(\ringosc.dstage[0].id.d0 ),
    .TE(\itrim[13] ),
    .Z(\ringosc.dstage[0].id.d1 ));
 sky130_fd_sc_hd__einvn_2 \ringosc.dstage[0].id.delayenb0  (.A(\ringosc.dstage[0].id.ts ),
    .TE_B(\itrim[0] ),
    .Z(\ringosc.dstage[0].id.out ));
 sky130_fd_sc_hd__einvn_1 \ringosc.dstage[0].id.delayenb1  (.A(\ringosc.dstage[0].id.ts ),
    .TE_B(\itrim[13] ),
    .Z(\ringosc.dstage[0].id.d1 ));
 sky130_fd_sc_hd__inv_1 \ringosc.dstage[0].id.delayint0  (.A(\ringosc.dstage[0].id.d1 ),
    .Y(\ringosc.dstage[0].id.d2 ));
 sky130_fd_sc_hd__clkbuf_1 \ringosc.dstage[10].id.delaybuf0  (.A(\ringosc.dstage[10].id.in ),
    .X(\ringosc.dstage[10].id.ts ));
 sky130_fd_sc_hd__clkbuf_1 \ringosc.dstage[10].id.delaybuf1  (.A(\ringosc.dstage[10].id.ts ),
    .X(\ringosc.dstage[10].id.d0 ));
 sky130_fd_sc_hd__einvp_2 \ringosc.dstage[10].id.delayen0  (.A(\ringosc.dstage[10].id.d2 ),
    .TE(\itrim[10] ),
    .Z(\ringosc.dstage[10].id.out ));
 sky130_fd_sc_hd__einvp_1 \ringosc.dstage[10].id.delayen1  (.A(\ringosc.dstage[10].id.d0 ),
    .TE(\itrim[23] ),
    .Z(\ringosc.dstage[10].id.d1 ));
 sky130_fd_sc_hd__einvn_2 \ringosc.dstage[10].id.delayenb0  (.A(\ringosc.dstage[10].id.ts ),
    .TE_B(\itrim[10] ),
    .Z(\ringosc.dstage[10].id.out ));
 sky130_fd_sc_hd__einvn_1 \ringosc.dstage[10].id.delayenb1  (.A(\ringosc.dstage[10].id.ts ),
    .TE_B(\itrim[23] ),
    .Z(\ringosc.dstage[10].id.d1 ));
 sky130_fd_sc_hd__inv_1 \ringosc.dstage[10].id.delayint0  (.A(\ringosc.dstage[10].id.d1 ),
    .Y(\ringosc.dstage[10].id.d2 ));
 sky130_fd_sc_hd__clkbuf_2 \ringosc.dstage[11].id.delaybuf0  (.A(\ringosc.dstage[10].id.out ),
    .X(\ringosc.dstage[11].id.ts ));
 sky130_fd_sc_hd__clkbuf_1 \ringosc.dstage[11].id.delaybuf1  (.A(\ringosc.dstage[11].id.ts ),
    .X(\ringosc.dstage[11].id.d0 ));
 sky130_fd_sc_hd__einvp_8 \ringosc.dstage[11].id.delayen0  (.A(\ringosc.dstage[11].id.d2 ),
    .TE(\itrim[11] ),
    .Z(\ringosc.dstage[11].id.out ));
 sky130_fd_sc_hd__einvp_1 \ringosc.dstage[11].id.delayen1  (.A(\ringosc.dstage[11].id.d0 ),
    .TE(\itrim[24] ),
    .Z(\ringosc.dstage[11].id.d1 ));
 sky130_fd_sc_hd__einvn_8 \ringosc.dstage[11].id.delayenb0  (.A(\ringosc.dstage[11].id.ts ),
    .TE_B(\itrim[11] ),
    .Z(\ringosc.dstage[11].id.out ));
 sky130_fd_sc_hd__einvn_1 \ringosc.dstage[11].id.delayenb1  (.A(\ringosc.dstage[11].id.ts ),
    .TE_B(\itrim[24] ),
    .Z(\ringosc.dstage[11].id.d1 ));
 sky130_fd_sc_hd__clkinv_1 \ringosc.dstage[11].id.delayint0  (.A(\ringosc.dstage[11].id.d1 ),
    .Y(\ringosc.dstage[11].id.d2 ));
 sky130_fd_sc_hd__clkbuf_1 \ringosc.dstage[1].id.delaybuf0  (.A(\ringosc.dstage[0].id.out ),
    .X(\ringosc.dstage[1].id.ts ));
 sky130_fd_sc_hd__clkbuf_1 \ringosc.dstage[1].id.delaybuf1  (.A(\ringosc.dstage[1].id.ts ),
    .X(\ringosc.dstage[1].id.d0 ));
 sky130_fd_sc_hd__einvp_2 \ringosc.dstage[1].id.delayen0  (.A(\ringosc.dstage[1].id.d2 ),
    .TE(\itrim[1] ),
    .Z(\ringosc.dstage[1].id.out ));
 sky130_fd_sc_hd__einvp_1 \ringosc.dstage[1].id.delayen1  (.A(\ringosc.dstage[1].id.d0 ),
    .TE(\itrim[14] ),
    .Z(\ringosc.dstage[1].id.d1 ));
 sky130_fd_sc_hd__einvn_2 \ringosc.dstage[1].id.delayenb0  (.A(\ringosc.dstage[1].id.ts ),
    .TE_B(\itrim[1] ),
    .Z(\ringosc.dstage[1].id.out ));
 sky130_fd_sc_hd__einvn_1 \ringosc.dstage[1].id.delayenb1  (.A(\ringosc.dstage[1].id.ts ),
    .TE_B(\itrim[14] ),
    .Z(\ringosc.dstage[1].id.d1 ));
 sky130_fd_sc_hd__inv_1 \ringosc.dstage[1].id.delayint0  (.A(\ringosc.dstage[1].id.d1 ),
    .Y(\ringosc.dstage[1].id.d2 ));
 sky130_fd_sc_hd__clkbuf_1 \ringosc.dstage[2].id.delaybuf0  (.A(\ringosc.dstage[1].id.out ),
    .X(\ringosc.dstage[2].id.ts ));
 sky130_fd_sc_hd__clkbuf_1 \ringosc.dstage[2].id.delaybuf1  (.A(\ringosc.dstage[2].id.ts ),
    .X(\ringosc.dstage[2].id.d0 ));
 sky130_fd_sc_hd__einvp_2 \ringosc.dstage[2].id.delayen0  (.A(\ringosc.dstage[2].id.d2 ),
    .TE(\itrim[2] ),
    .Z(\ringosc.dstage[2].id.out ));
 sky130_fd_sc_hd__einvp_1 \ringosc.dstage[2].id.delayen1  (.A(\ringosc.dstage[2].id.d0 ),
    .TE(\itrim[15] ),
    .Z(\ringosc.dstage[2].id.d1 ));
 sky130_fd_sc_hd__einvn_2 \ringosc.dstage[2].id.delayenb0  (.A(\ringosc.dstage[2].id.ts ),
    .TE_B(\itrim[2] ),
    .Z(\ringosc.dstage[2].id.out ));
 sky130_fd_sc_hd__einvn_1 \ringosc.dstage[2].id.delayenb1  (.A(\ringosc.dstage[2].id.ts ),
    .TE_B(\itrim[15] ),
    .Z(\ringosc.dstage[2].id.d1 ));
 sky130_fd_sc_hd__inv_1 \ringosc.dstage[2].id.delayint0  (.A(\ringosc.dstage[2].id.d1 ),
    .Y(\ringosc.dstage[2].id.d2 ));
 sky130_fd_sc_hd__clkbuf_1 \ringosc.dstage[3].id.delaybuf0  (.A(\ringosc.dstage[2].id.out ),
    .X(\ringosc.dstage[3].id.ts ));
 sky130_fd_sc_hd__clkbuf_1 \ringosc.dstage[3].id.delaybuf1  (.A(\ringosc.dstage[3].id.ts ),
    .X(\ringosc.dstage[3].id.d0 ));
 sky130_fd_sc_hd__einvp_2 \ringosc.dstage[3].id.delayen0  (.A(\ringosc.dstage[3].id.d2 ),
    .TE(\itrim[3] ),
    .Z(\ringosc.dstage[3].id.out ));
 sky130_fd_sc_hd__einvp_1 \ringosc.dstage[3].id.delayen1  (.A(\ringosc.dstage[3].id.d0 ),
    .TE(\itrim[16] ),
    .Z(\ringosc.dstage[3].id.d1 ));
 sky130_fd_sc_hd__einvn_2 \ringosc.dstage[3].id.delayenb0  (.A(\ringosc.dstage[3].id.ts ),
    .TE_B(\itrim[3] ),
    .Z(\ringosc.dstage[3].id.out ));
 sky130_fd_sc_hd__einvn_1 \ringosc.dstage[3].id.delayenb1  (.A(\ringosc.dstage[3].id.ts ),
    .TE_B(\itrim[16] ),
    .Z(\ringosc.dstage[3].id.d1 ));
 sky130_fd_sc_hd__inv_1 \ringosc.dstage[3].id.delayint0  (.A(\ringosc.dstage[3].id.d1 ),
    .Y(\ringosc.dstage[3].id.d2 ));
 sky130_fd_sc_hd__clkbuf_1 \ringosc.dstage[4].id.delaybuf0  (.A(\ringosc.dstage[3].id.out ),
    .X(\ringosc.dstage[4].id.ts ));
 sky130_fd_sc_hd__clkbuf_1 \ringosc.dstage[4].id.delaybuf1  (.A(\ringosc.dstage[4].id.ts ),
    .X(\ringosc.dstage[4].id.d0 ));
 sky130_fd_sc_hd__einvp_2 \ringosc.dstage[4].id.delayen0  (.A(\ringosc.dstage[4].id.d2 ),
    .TE(\itrim[4] ),
    .Z(\ringosc.dstage[4].id.out ));
 sky130_fd_sc_hd__einvp_1 \ringosc.dstage[4].id.delayen1  (.A(\ringosc.dstage[4].id.d0 ),
    .TE(\itrim[17] ),
    .Z(\ringosc.dstage[4].id.d1 ));
 sky130_fd_sc_hd__einvn_2 \ringosc.dstage[4].id.delayenb0  (.A(\ringosc.dstage[4].id.ts ),
    .TE_B(\itrim[4] ),
    .Z(\ringosc.dstage[4].id.out ));
 sky130_fd_sc_hd__einvn_1 \ringosc.dstage[4].id.delayenb1  (.A(\ringosc.dstage[4].id.ts ),
    .TE_B(\itrim[17] ),
    .Z(\ringosc.dstage[4].id.d1 ));
 sky130_fd_sc_hd__inv_1 \ringosc.dstage[4].id.delayint0  (.A(\ringosc.dstage[4].id.d1 ),
    .Y(\ringosc.dstage[4].id.d2 ));
 sky130_fd_sc_hd__clkbuf_1 \ringosc.dstage[5].id.delaybuf0  (.A(\ringosc.dstage[4].id.out ),
    .X(\ringosc.dstage[5].id.ts ));
 sky130_fd_sc_hd__clkbuf_1 \ringosc.dstage[5].id.delaybuf1  (.A(\ringosc.dstage[5].id.ts ),
    .X(\ringosc.dstage[5].id.d0 ));
 sky130_fd_sc_hd__einvp_2 \ringosc.dstage[5].id.delayen0  (.A(\ringosc.dstage[5].id.d2 ),
    .TE(\itrim[5] ),
    .Z(\ringosc.dstage[5].id.out ));
 sky130_fd_sc_hd__einvp_1 \ringosc.dstage[5].id.delayen1  (.A(\ringosc.dstage[5].id.d0 ),
    .TE(\itrim[18] ),
    .Z(\ringosc.dstage[5].id.d1 ));
 sky130_fd_sc_hd__einvn_2 \ringosc.dstage[5].id.delayenb0  (.A(\ringosc.dstage[5].id.ts ),
    .TE_B(\itrim[5] ),
    .Z(\ringosc.dstage[5].id.out ));
 sky130_fd_sc_hd__einvn_1 \ringosc.dstage[5].id.delayenb1  (.A(\ringosc.dstage[5].id.ts ),
    .TE_B(\itrim[18] ),
    .Z(\ringosc.dstage[5].id.d1 ));
 sky130_fd_sc_hd__inv_1 \ringosc.dstage[5].id.delayint0  (.A(\ringosc.dstage[5].id.d1 ),
    .Y(\ringosc.dstage[5].id.d2 ));
 sky130_fd_sc_hd__clkbuf_1 \ringosc.dstage[6].id.delaybuf0  (.A(\ringosc.dstage[5].id.out ),
    .X(\ringosc.dstage[6].id.ts ));
 sky130_fd_sc_hd__clkbuf_1 \ringosc.dstage[6].id.delaybuf1  (.A(\ringosc.dstage[6].id.ts ),
    .X(\ringosc.dstage[6].id.d0 ));
 sky130_fd_sc_hd__einvp_2 \ringosc.dstage[6].id.delayen0  (.A(\ringosc.dstage[6].id.d2 ),
    .TE(\itrim[6] ),
    .Z(\ringosc.dstage[6].id.out ));
 sky130_fd_sc_hd__einvp_1 \ringosc.dstage[6].id.delayen1  (.A(\ringosc.dstage[6].id.d0 ),
    .TE(\itrim[19] ),
    .Z(\ringosc.dstage[6].id.d1 ));
 sky130_fd_sc_hd__einvn_2 \ringosc.dstage[6].id.delayenb0  (.A(\ringosc.dstage[6].id.ts ),
    .TE_B(\itrim[6] ),
    .Z(\ringosc.dstage[6].id.out ));
 sky130_fd_sc_hd__einvn_1 \ringosc.dstage[6].id.delayenb1  (.A(\ringosc.dstage[6].id.ts ),
    .TE_B(\itrim[19] ),
    .Z(\ringosc.dstage[6].id.d1 ));
 sky130_fd_sc_hd__inv_1 \ringosc.dstage[6].id.delayint0  (.A(\ringosc.dstage[6].id.d1 ),
    .Y(\ringosc.dstage[6].id.d2 ));
 sky130_fd_sc_hd__clkbuf_1 \ringosc.dstage[7].id.delaybuf0  (.A(\ringosc.dstage[6].id.out ),
    .X(\ringosc.dstage[7].id.ts ));
 sky130_fd_sc_hd__clkbuf_1 \ringosc.dstage[7].id.delaybuf1  (.A(\ringosc.dstage[7].id.ts ),
    .X(\ringosc.dstage[7].id.d0 ));
 sky130_fd_sc_hd__einvp_2 \ringosc.dstage[7].id.delayen0  (.A(\ringosc.dstage[7].id.d2 ),
    .TE(\itrim[7] ),
    .Z(\ringosc.dstage[7].id.out ));
 sky130_fd_sc_hd__einvp_1 \ringosc.dstage[7].id.delayen1  (.A(\ringosc.dstage[7].id.d0 ),
    .TE(\itrim[20] ),
    .Z(\ringosc.dstage[7].id.d1 ));
 sky130_fd_sc_hd__einvn_2 \ringosc.dstage[7].id.delayenb0  (.A(\ringosc.dstage[7].id.ts ),
    .TE_B(\itrim[7] ),
    .Z(\ringosc.dstage[7].id.out ));
 sky130_fd_sc_hd__einvn_1 \ringosc.dstage[7].id.delayenb1  (.A(\ringosc.dstage[7].id.ts ),
    .TE_B(\itrim[20] ),
    .Z(\ringosc.dstage[7].id.d1 ));
 sky130_fd_sc_hd__inv_1 \ringosc.dstage[7].id.delayint0  (.A(\ringosc.dstage[7].id.d1 ),
    .Y(\ringosc.dstage[7].id.d2 ));
 sky130_fd_sc_hd__clkbuf_1 \ringosc.dstage[8].id.delaybuf0  (.A(\ringosc.dstage[7].id.out ),
    .X(\ringosc.dstage[8].id.ts ));
 sky130_fd_sc_hd__clkbuf_1 \ringosc.dstage[8].id.delaybuf1  (.A(\ringosc.dstage[8].id.ts ),
    .X(\ringosc.dstage[8].id.d0 ));
 sky130_fd_sc_hd__einvp_2 \ringosc.dstage[8].id.delayen0  (.A(\ringosc.dstage[8].id.d2 ),
    .TE(\itrim[8] ),
    .Z(\ringosc.dstage[8].id.out ));
 sky130_fd_sc_hd__einvp_1 \ringosc.dstage[8].id.delayen1  (.A(\ringosc.dstage[8].id.d0 ),
    .TE(\itrim[21] ),
    .Z(\ringosc.dstage[8].id.d1 ));
 sky130_fd_sc_hd__einvn_2 \ringosc.dstage[8].id.delayenb0  (.A(\ringosc.dstage[8].id.ts ),
    .TE_B(\itrim[8] ),
    .Z(\ringosc.dstage[8].id.out ));
 sky130_fd_sc_hd__einvn_1 \ringosc.dstage[8].id.delayenb1  (.A(\ringosc.dstage[8].id.ts ),
    .TE_B(\itrim[21] ),
    .Z(\ringosc.dstage[8].id.d1 ));
 sky130_fd_sc_hd__inv_1 \ringosc.dstage[8].id.delayint0  (.A(\ringosc.dstage[8].id.d1 ),
    .Y(\ringosc.dstage[8].id.d2 ));
 sky130_fd_sc_hd__clkbuf_1 \ringosc.dstage[9].id.delaybuf0  (.A(\ringosc.dstage[8].id.out ),
    .X(\ringosc.dstage[9].id.ts ));
 sky130_fd_sc_hd__clkbuf_1 \ringosc.dstage[9].id.delaybuf1  (.A(\ringosc.dstage[9].id.ts ),
    .X(\ringosc.dstage[9].id.d0 ));
 sky130_fd_sc_hd__einvp_2 \ringosc.dstage[9].id.delayen0  (.A(\ringosc.dstage[9].id.d2 ),
    .TE(\itrim[9] ),
    .Z(\ringosc.dstage[10].id.in ));
 sky130_fd_sc_hd__einvp_1 \ringosc.dstage[9].id.delayen1  (.A(\ringosc.dstage[9].id.d0 ),
    .TE(\itrim[22] ),
    .Z(\ringosc.dstage[9].id.d1 ));
 sky130_fd_sc_hd__einvn_2 \ringosc.dstage[9].id.delayenb0  (.A(\ringosc.dstage[9].id.ts ),
    .TE_B(\itrim[9] ),
    .Z(\ringosc.dstage[10].id.in ));
 sky130_fd_sc_hd__einvn_1 \ringosc.dstage[9].id.delayenb1  (.A(\ringosc.dstage[9].id.ts ),
    .TE_B(\itrim[22] ),
    .Z(\ringosc.dstage[9].id.d1 ));
 sky130_fd_sc_hd__inv_1 \ringosc.dstage[9].id.delayint0  (.A(\ringosc.dstage[9].id.d1 ),
    .Y(\ringosc.dstage[9].id.d2 ));
 sky130_fd_sc_hd__clkinv_2 \ringosc.ibufp00  (.A(\ringosc.dstage[0].id.in ),
    .Y(\ringosc.c[0] ));
 sky130_fd_sc_hd__clkinv_8 \ringosc.ibufp01  (.A(\ringosc.c[0] ),
    .Y(\clockp_buffer_in[0] ));
 sky130_fd_sc_hd__clkinv_2 \ringosc.ibufp10  (.A(\ringosc.dstage[5].id.out ),
    .Y(\ringosc.c[1] ));
 sky130_fd_sc_hd__clkinv_4 \ringosc.ibufp11  (.A(\ringosc.c[1] ),
    .Y(\clockp_buffer_in[1] ));
 sky130_fd_sc_hd__conb_1 \ringosc.iss.const1  (.HI(\ringosc.iss.one ));
 sky130_fd_sc_hd__or2_1 \ringosc.iss.ctrlen0  (.A(net114),
    .B(\itrim[12] ),
    .X(\ringosc.iss.ctrl0 ));
 sky130_fd_sc_hd__clkbuf_1 \ringosc.iss.delaybuf0  (.A(\ringosc.dstage[11].id.out ),
    .X(\ringosc.iss.d0 ));
 sky130_fd_sc_hd__einvp_4 \ringosc.iss.delayen0  (.A(\ringosc.iss.d2 ),
    .TE(\itrim[12] ),
    .Z(\ringosc.dstage[0].id.in ));
 sky130_fd_sc_hd__einvp_1 \ringosc.iss.delayen1  (.A(\ringosc.iss.d0 ),
    .TE(\itrim[25] ),
    .Z(\ringosc.iss.d1 ));
 sky130_fd_sc_hd__einvn_4 \ringosc.iss.delayenb0  (.A(\ringosc.dstage[11].id.out ),
    .TE_B(\ringosc.iss.ctrl0 ),
    .Z(\ringosc.dstage[0].id.in ));
 sky130_fd_sc_hd__einvn_1 \ringosc.iss.delayenb1  (.A(\ringosc.dstage[11].id.out ),
    .TE_B(\itrim[25] ),
    .Z(\ringosc.iss.d1 ));
 sky130_fd_sc_hd__inv_1 \ringosc.iss.delayint0  (.A(\ringosc.iss.d1 ),
    .Y(\ringosc.iss.d2 ));
 sky130_fd_sc_hd__einvp_4 \ringosc.iss.reseten0  (.A(\ringosc.iss.one ),
    .TE(net114),
    .Z(\ringosc.dstage[0].id.in ));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_242 ();
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout104 (.A(net106),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_1 fanout105 (.A(net106),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_1 fanout106 (.A(net107),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_1 fanout107 (.A(\dll_control.tint[4] ),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_2 fanout108 (.A(net109),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_1 fanout109 (.A(\dll_control.tint[3] ),
    .X(net109));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout110 (.A(\dll_control.tint[2] ),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_2 fanout111 (.A(\dll_control.tint[1] ),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_1 fanout112 (.A(\dll_control.tint[1] ),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_2 fanout113 (.A(\dll_control.tint[0] ),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_2 fanout114 (.A(ireset),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_2 fanout115 (.A(net116),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_2 fanout116 (.A(net125),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_1 fanout117 (.A(net125),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_2 fanout118 (.A(net124),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_1 fanout119 (.A(net124),
    .X(net119));
 sky130_fd_sc_hd__clkbuf_2 fanout120 (.A(net121),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_1 fanout121 (.A(net122),
    .X(net121));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout122 (.A(net123),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_1 fanout123 (.A(net124),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_1 fanout124 (.A(net125),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_1 fanout125 (.A(dco),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_2 fanout126 (.A(net129),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_2 fanout127 (.A(net128),
    .X(net127));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout128 (.A(net129),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_1 fanout129 (.A(net139),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_2 fanout130 (.A(net134),
    .X(net130));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout131 (.A(net134),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_2 fanout132 (.A(net133),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_2 fanout133 (.A(net134),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_1 fanout134 (.A(net139),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_2 fanout135 (.A(net136),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_1 fanout136 (.A(net138),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_2 fanout137 (.A(net138),
    .X(net137));
 sky130_fd_sc_hd__clkbuf_1 fanout138 (.A(net139),
    .X(net138));
 sky130_fd_sc_hd__clkbuf_1 fanout139 (.A(dco),
    .X(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(enable));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(ext_trim[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(ext_trim[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(ext_trim[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(ext_trim[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(ext_trim[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(ext_trim[25]));
 sky130_fd_sc_hd__fill_1 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_107 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_14 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_140 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_247 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_140 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_265 ();
endmodule
