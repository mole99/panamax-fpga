magic
tech sky130A
magscale 1 2
timestamp 1746622459
<< viali >>
rect 5549 20553 5583 20587
rect 8677 20553 8711 20587
rect 10103 20553 10137 20587
rect 12081 20553 12115 20587
rect 14197 20553 14231 20587
rect 16129 20553 16163 20587
rect 12725 20485 12759 20519
rect 4445 20417 4479 20451
rect 5549 20417 5583 20451
rect 6009 20417 6043 20451
rect 6586 20417 6620 20451
rect 7389 20417 7423 20451
rect 7941 20417 7975 20451
rect 9137 20417 9171 20451
rect 9714 20417 9748 20451
rect 10174 20417 10208 20451
rect 14841 20417 14875 20451
rect 15434 20417 15468 20451
rect 4629 20349 4663 20383
rect 5181 20349 5215 20383
rect 8309 20349 8343 20383
rect 11713 20349 11747 20383
rect 12357 20349 12391 20383
rect 14565 20349 14599 20383
rect 15761 20349 15795 20383
rect 8677 20281 8711 20315
rect 12081 20281 12115 20315
rect 14197 20281 14231 20315
rect 16129 20281 16163 20315
rect 5365 20213 5399 20247
rect 5825 20213 5859 20247
rect 6515 20213 6549 20247
rect 7389 20213 7423 20247
rect 9321 20213 9355 20247
rect 9643 20213 9677 20247
rect 12725 20213 12759 20247
rect 15025 20213 15059 20247
rect 15347 20213 15381 20247
rect 6193 20009 6227 20043
rect 9873 20009 9907 20043
rect 12173 20009 12207 20043
rect 14197 20009 14231 20043
rect 15485 20009 15519 20043
rect 16313 20009 16347 20043
rect 17233 20009 17267 20043
rect 4813 19941 4847 19975
rect 5549 19941 5583 19975
rect 7757 19941 7791 19975
rect 8493 19941 8527 19975
rect 9413 19941 9447 19975
rect 10333 19941 10367 19975
rect 11161 19941 11195 19975
rect 12449 19941 12483 19975
rect 13737 19941 13771 19975
rect 16497 19941 16531 19975
rect 5641 19873 5675 19907
rect 7573 19873 7607 19907
rect 8033 19873 8067 19907
rect 8585 19873 8619 19907
rect 10057 19873 10091 19907
rect 15209 19873 15243 19907
rect 15485 19873 15519 19907
rect 15853 19873 15887 19907
rect 4261 19805 4295 19839
rect 4813 19805 4847 19839
rect 5089 19805 5123 19839
rect 5549 19805 5583 19839
rect 6009 19805 6043 19839
rect 6745 19805 6779 19839
rect 7205 19805 7239 19839
rect 7757 19805 7791 19839
rect 9045 19805 9079 19839
rect 9689 19805 9723 19839
rect 10517 19805 10551 19839
rect 11345 19805 11379 19839
rect 11713 19805 11747 19839
rect 11989 19805 12023 19839
rect 12449 19805 12483 19839
rect 13001 19805 13035 19839
rect 13277 19805 13311 19839
rect 14381 19805 14415 19839
rect 14657 19805 14691 19839
rect 16129 19805 16163 19839
rect 16890 19805 16924 19839
rect 17417 19805 17451 19839
rect 11437 19737 11471 19771
rect 11529 19737 11563 19771
rect 13829 19737 13863 19771
rect 15117 19737 15151 19771
rect 16497 19737 16531 19771
rect 6929 19669 6963 19703
rect 9413 19669 9447 19703
rect 16819 19669 16853 19703
rect 5365 19465 5399 19499
rect 5733 19465 5767 19499
rect 7021 19465 7055 19499
rect 9965 19465 9999 19499
rect 11253 19465 11287 19499
rect 12265 19465 12299 19499
rect 13139 19465 13173 19499
rect 16405 19465 16439 19499
rect 4445 19397 4479 19431
rect 7757 19397 7791 19431
rect 9229 19397 9263 19431
rect 10767 19397 10801 19431
rect 10977 19397 11011 19431
rect 11779 19397 11813 19431
rect 12541 19397 12575 19431
rect 14657 19397 14691 19431
rect 16773 19397 16807 19431
rect 4353 19329 4387 19363
rect 5825 19329 5859 19363
rect 6837 19329 6871 19363
rect 7481 19329 7515 19363
rect 7849 19329 7883 19363
rect 8309 19329 8343 19363
rect 9045 19329 9079 19363
rect 9321 19329 9355 19363
rect 10885 19329 10919 19363
rect 11069 19329 11103 19363
rect 11897 19329 11931 19363
rect 11989 19329 12023 19363
rect 12081 19329 12115 19363
rect 13036 19329 13070 19363
rect 14197 19329 14231 19363
rect 14749 19329 14783 19363
rect 15393 19351 15427 19385
rect 15945 19329 15979 19363
rect 16221 19329 16255 19363
rect 17325 19329 17359 19363
rect 4997 19261 5031 19295
rect 5365 19261 5399 19295
rect 8861 19261 8895 19295
rect 9597 19261 9631 19295
rect 9965 19261 9999 19295
rect 10609 19261 10643 19295
rect 11621 19261 11655 19295
rect 15945 19193 15979 19227
rect 16865 19193 16899 19227
rect 7297 19125 7331 19159
rect 12633 19125 12667 19159
rect 4813 18921 4847 18955
rect 5457 18921 5491 18955
rect 5733 18921 5767 18955
rect 7113 18921 7147 18955
rect 8585 18921 8619 18955
rect 9045 18921 9079 18955
rect 9413 18921 9447 18955
rect 10425 18921 10459 18955
rect 10609 18921 10643 18955
rect 12725 18921 12759 18955
rect 14749 18921 14783 18955
rect 10057 18853 10091 18887
rect 7757 18785 7791 18819
rect 9505 18785 9539 18819
rect 10977 18785 11011 18819
rect 3376 18717 3410 18751
rect 4445 18717 4479 18751
rect 4813 18717 4847 18751
rect 5273 18717 5307 18751
rect 5733 18717 5767 18751
rect 5917 18717 5951 18751
rect 8125 18717 8159 18751
rect 8217 18717 8251 18751
rect 8401 18717 8435 18751
rect 9229 18717 9263 18751
rect 11253 18717 11287 18751
rect 11529 18717 11563 18751
rect 11713 18717 11747 18751
rect 12173 18717 12207 18751
rect 12357 18717 12391 18751
rect 12449 18717 12483 18751
rect 12541 18717 12575 18751
rect 13001 18717 13035 18751
rect 13185 18717 13219 18751
rect 14197 18717 14231 18751
rect 14565 18717 14599 18751
rect 16773 18717 16807 18751
rect 17417 18717 17451 18751
rect 17728 18717 17762 18751
rect 3479 18649 3513 18683
rect 3893 18649 3927 18683
rect 3985 18649 4019 18683
rect 7481 18649 7515 18683
rect 10425 18649 10459 18683
rect 11411 18649 11445 18683
rect 11621 18649 11655 18683
rect 11897 18649 11931 18683
rect 13093 18649 13127 18683
rect 14381 18649 14415 18683
rect 14473 18649 14507 18683
rect 15025 18649 15059 18683
rect 15209 18649 15243 18683
rect 6745 18581 6779 18615
rect 7573 18581 7607 18615
rect 10609 18581 10643 18615
rect 16957 18581 16991 18615
rect 17233 18581 17267 18615
rect 17831 18581 17865 18615
rect 3249 18377 3283 18411
rect 5457 18377 5491 18411
rect 6469 18377 6503 18411
rect 11043 18377 11077 18411
rect 12265 18377 12299 18411
rect 12541 18377 12575 18411
rect 13093 18377 13127 18411
rect 14197 18377 14231 18411
rect 15301 18377 15335 18411
rect 3985 18309 4019 18343
rect 4445 18309 4479 18343
rect 11253 18309 11287 18343
rect 13369 18309 13403 18343
rect 16405 18309 16439 18343
rect 18153 18309 18187 18343
rect 3249 18241 3283 18275
rect 3525 18241 3559 18275
rect 4077 18241 4111 18275
rect 4353 18241 4387 18275
rect 4629 18241 4663 18275
rect 5917 18241 5951 18275
rect 6837 18241 6871 18275
rect 7481 18241 7515 18275
rect 8953 18241 8987 18275
rect 9413 18241 9447 18275
rect 9597 18241 9631 18275
rect 10241 18241 10275 18275
rect 10425 18241 10459 18275
rect 11621 18241 11655 18275
rect 11805 18241 11839 18275
rect 11897 18241 11931 18275
rect 12035 18241 12069 18275
rect 12541 18241 12575 18275
rect 12633 18241 12667 18275
rect 12817 18241 12851 18275
rect 13231 18241 13265 18275
rect 13461 18241 13495 18275
rect 13644 18241 13678 18275
rect 13737 18241 13771 18275
rect 14013 18241 14047 18275
rect 14473 18241 14507 18275
rect 14565 18241 14599 18275
rect 14749 18241 14783 18275
rect 15209 18241 15243 18275
rect 15485 18241 15519 18275
rect 15669 18241 15703 18275
rect 16773 18241 16807 18275
rect 17325 18241 17359 18275
rect 2881 18173 2915 18207
rect 4813 18173 4847 18207
rect 5089 18173 5123 18207
rect 6929 18173 6963 18207
rect 7021 18173 7055 18207
rect 9781 18173 9815 18207
rect 14933 18173 14967 18207
rect 16037 18173 16071 18207
rect 17601 18173 17635 18207
rect 3249 18105 3283 18139
rect 5457 18105 5491 18139
rect 5733 18105 5767 18139
rect 9137 18105 9171 18139
rect 10885 18105 10919 18139
rect 17325 18105 17359 18139
rect 18061 18105 18095 18139
rect 10609 18037 10643 18071
rect 11069 18037 11103 18071
rect 12725 18037 12759 18071
rect 16405 18037 16439 18071
rect 5365 17833 5399 17867
rect 9045 17833 9079 17867
rect 9965 17833 9999 17867
rect 11529 17833 11563 17867
rect 11989 17833 12023 17867
rect 13737 17833 13771 17867
rect 15393 17833 15427 17867
rect 15945 17833 15979 17867
rect 4261 17765 4295 17799
rect 7573 17765 7607 17799
rect 8493 17765 8527 17799
rect 9781 17765 9815 17799
rect 12541 17765 12575 17799
rect 17049 17765 17083 17799
rect 4077 17697 4111 17731
rect 7849 17697 7883 17731
rect 10517 17697 10551 17731
rect 15945 17697 15979 17731
rect 16681 17697 16715 17731
rect 4445 17629 4479 17663
rect 4838 17629 4872 17663
rect 5181 17629 5215 17663
rect 5641 17629 5675 17663
rect 5733 17629 5767 17663
rect 5917 17629 5951 17663
rect 6929 17629 6963 17663
rect 7205 17629 7239 17663
rect 8217 17629 8251 17663
rect 8677 17629 8711 17663
rect 9229 17629 9263 17663
rect 9413 17629 9447 17663
rect 9505 17629 9539 17663
rect 10425 17629 10459 17663
rect 10609 17629 10643 17663
rect 10885 17629 10919 17663
rect 11069 17629 11103 17663
rect 12173 17629 12207 17663
rect 12265 17629 12299 17663
rect 12817 17629 12851 17663
rect 13001 17629 13035 17663
rect 13461 17629 13495 17663
rect 14197 17629 14231 17663
rect 14290 17629 14324 17663
rect 14662 17629 14696 17663
rect 15577 17629 15611 17663
rect 16129 17629 16163 17663
rect 16405 17629 16439 17663
rect 17969 17629 18003 17663
rect 18613 17629 18647 17663
rect 9919 17595 9953 17629
rect 10149 17561 10183 17595
rect 11345 17561 11379 17595
rect 11561 17561 11595 17595
rect 13737 17561 13771 17595
rect 14473 17561 14507 17595
rect 14565 17561 14599 17595
rect 18153 17561 18187 17595
rect 4767 17493 4801 17527
rect 6101 17493 6135 17527
rect 6745 17493 6779 17527
rect 7573 17493 7607 17527
rect 7849 17493 7883 17527
rect 10885 17493 10919 17527
rect 11713 17493 11747 17527
rect 12173 17493 12207 17527
rect 12357 17493 12391 17527
rect 12909 17493 12943 17527
rect 13553 17493 13587 17527
rect 14841 17493 14875 17527
rect 16313 17493 16347 17527
rect 17049 17493 17083 17527
rect 18429 17493 18463 17527
rect 4721 17289 4755 17323
rect 8861 17289 8895 17323
rect 11989 17289 12023 17323
rect 12541 17289 12575 17323
rect 3525 17221 3559 17255
rect 4353 17221 4387 17255
rect 4445 17221 4479 17255
rect 7021 17221 7055 17255
rect 14289 17221 14323 17255
rect 3065 17153 3099 17187
rect 3617 17153 3651 17187
rect 5089 17153 5123 17187
rect 5365 17153 5399 17187
rect 5917 17153 5951 17187
rect 6520 17153 6554 17187
rect 7941 17153 7975 17187
rect 8125 17153 8159 17187
rect 8401 17153 8435 17187
rect 8585 17153 8619 17187
rect 9045 17153 9079 17187
rect 9137 17153 9171 17187
rect 9229 17153 9263 17187
rect 9413 17153 9447 17187
rect 9689 17153 9723 17187
rect 9873 17153 9907 17187
rect 9965 17153 9999 17187
rect 10057 17153 10091 17187
rect 10609 17153 10643 17187
rect 11069 17153 11103 17187
rect 11897 17153 11931 17187
rect 12725 17153 12759 17187
rect 12817 17153 12851 17187
rect 12909 17153 12943 17187
rect 13461 17153 13495 17187
rect 13553 17153 13587 17187
rect 14013 17153 14047 17187
rect 14197 17153 14231 17187
rect 14381 17153 14415 17187
rect 16922 17153 16956 17187
rect 17325 17153 17359 17187
rect 18245 17153 18279 17187
rect 19349 17153 19383 17187
rect 20729 17153 20763 17187
rect 3893 17085 3927 17119
rect 4721 17085 4755 17119
rect 6607 17085 6641 17119
rect 6929 17085 6963 17119
rect 7481 17085 7515 17119
rect 8033 17085 8067 17119
rect 11780 17085 11814 17119
rect 12265 17085 12299 17119
rect 13277 17085 13311 17119
rect 18889 17085 18923 17119
rect 19257 17085 19291 17119
rect 10241 17017 10275 17051
rect 11161 17017 11195 17051
rect 11621 17017 11655 17051
rect 13369 17017 13403 17051
rect 18613 17017 18647 17051
rect 5917 16949 5951 16983
rect 8493 16949 8527 16983
rect 10701 16949 10735 16983
rect 14565 16949 14599 16983
rect 16819 16949 16853 16983
rect 4445 16745 4479 16779
rect 4813 16745 4847 16779
rect 7113 16745 7147 16779
rect 9597 16745 9631 16779
rect 11161 16745 11195 16779
rect 11621 16745 11655 16779
rect 5273 16677 5307 16711
rect 6193 16677 6227 16711
rect 10609 16677 10643 16711
rect 13461 16677 13495 16711
rect 14473 16677 14507 16711
rect 16497 16677 16531 16711
rect 16957 16677 16991 16711
rect 18429 16677 18463 16711
rect 7849 16609 7883 16643
rect 16773 16609 16807 16643
rect 17417 16609 17451 16643
rect 18061 16609 18095 16643
rect 3985 16541 4019 16575
rect 4261 16541 4295 16575
rect 4997 16541 5031 16575
rect 5457 16541 5491 16575
rect 5733 16541 5767 16575
rect 6561 16541 6595 16575
rect 7113 16541 7147 16575
rect 7389 16541 7423 16575
rect 7665 16541 7699 16575
rect 8493 16541 8527 16575
rect 8677 16541 8711 16575
rect 9045 16541 9079 16575
rect 9229 16541 9263 16575
rect 9413 16541 9447 16575
rect 9873 16541 9907 16575
rect 10149 16541 10183 16575
rect 10517 16541 10551 16575
rect 10701 16541 10735 16575
rect 11252 16541 11286 16575
rect 11345 16541 11379 16575
rect 11805 16541 11839 16575
rect 11989 16541 12023 16575
rect 12173 16541 12207 16575
rect 12724 16541 12758 16575
rect 12817 16541 12851 16575
rect 13093 16541 13127 16575
rect 13277 16541 13311 16575
rect 14749 16541 14783 16575
rect 15117 16541 15151 16575
rect 15945 16541 15979 16575
rect 16129 16541 16163 16575
rect 16221 16541 16255 16575
rect 16313 16541 16347 16575
rect 17785 16541 17819 16575
rect 18889 16541 18923 16575
rect 6285 16473 6319 16507
rect 7481 16473 7515 16507
rect 9321 16473 9355 16507
rect 11897 16473 11931 16507
rect 14933 16473 14967 16507
rect 15025 16473 15059 16507
rect 15669 16473 15703 16507
rect 17141 16473 17175 16507
rect 4077 16405 4111 16439
rect 8677 16405 8711 16439
rect 10149 16405 10183 16439
rect 12449 16405 12483 16439
rect 15301 16405 15335 16439
rect 17785 16405 17819 16439
rect 18429 16405 18463 16439
rect 18705 16405 18739 16439
rect 6101 16201 6135 16235
rect 6837 16201 6871 16235
rect 8769 16201 8803 16235
rect 10885 16201 10919 16235
rect 11621 16201 11655 16235
rect 13093 16201 13127 16235
rect 13369 16201 13403 16235
rect 14197 16201 14231 16235
rect 17141 16201 17175 16235
rect 9689 16133 9723 16167
rect 14841 16133 14875 16167
rect 16129 16133 16163 16167
rect 16405 16133 16439 16167
rect 3249 16065 3283 16099
rect 3433 16065 3467 16099
rect 4169 16065 4203 16099
rect 4353 16065 4387 16099
rect 6101 16065 6135 16099
rect 7297 16065 7331 16099
rect 7757 16065 7791 16099
rect 8953 16065 8987 16099
rect 9229 16065 9263 16099
rect 9413 16065 9447 16099
rect 9873 16065 9907 16099
rect 10149 16065 10183 16099
rect 11069 16065 11103 16099
rect 11253 16065 11287 16099
rect 11805 16065 11839 16099
rect 11897 16065 11931 16099
rect 12173 16065 12207 16099
rect 12633 16065 12667 16099
rect 12725 16065 12759 16099
rect 12817 16065 12851 16099
rect 14197 16065 14231 16099
rect 14381 16065 14415 16099
rect 15025 16065 15059 16099
rect 15209 16065 15243 16099
rect 15485 16065 15519 16099
rect 16773 16065 16807 16099
rect 17601 16065 17635 16099
rect 5733 15997 5767 16031
rect 6469 15997 6503 16031
rect 12081 15997 12115 16031
rect 12909 15997 12943 16031
rect 13829 15997 13863 16031
rect 6837 15929 6871 15963
rect 7113 15929 7147 15963
rect 7941 15929 7975 15963
rect 9965 15929 9999 15963
rect 10057 15929 10091 15963
rect 13461 15929 13495 15963
rect 17141 15929 17175 15963
rect 17417 15929 17451 15963
rect 3249 15861 3283 15895
rect 4353 15861 4387 15895
rect 6101 15861 6135 15895
rect 6423 15657 6457 15691
rect 8677 15657 8711 15691
rect 11161 15657 11195 15691
rect 12725 15657 12759 15691
rect 7021 15589 7055 15623
rect 9965 15589 9999 15623
rect 10517 15589 10551 15623
rect 12817 15589 12851 15623
rect 13461 15589 13495 15623
rect 3249 15521 3283 15555
rect 9597 15521 9631 15555
rect 10701 15521 10735 15555
rect 11437 15521 11471 15555
rect 14473 15521 14507 15555
rect 15577 15521 15611 15555
rect 16221 15521 16255 15555
rect 2513 15453 2547 15487
rect 2697 15453 2731 15487
rect 3157 15453 3191 15487
rect 3893 15453 3927 15487
rect 6494 15453 6528 15487
rect 8033 15453 8067 15487
rect 8217 15453 8251 15487
rect 8493 15453 8527 15487
rect 9137 15453 9171 15487
rect 9781 15453 9815 15487
rect 11069 15453 11103 15487
rect 11713 15453 11747 15487
rect 11897 15453 11931 15487
rect 12265 15453 12299 15487
rect 12357 15453 12391 15487
rect 13645 15453 13679 15487
rect 14197 15453 14231 15487
rect 16497 15453 16531 15487
rect 4169 15385 4203 15419
rect 7205 15385 7239 15419
rect 9321 15385 9355 15419
rect 10241 15385 10275 15419
rect 13185 15385 13219 15419
rect 2605 15317 2639 15351
rect 3525 15317 3559 15351
rect 5641 15317 5675 15351
rect 8125 15317 8159 15351
rect 11161 15317 11195 15351
rect 11253 15317 11287 15351
rect 8585 15113 8619 15147
rect 10057 15113 10091 15147
rect 11161 15113 11195 15147
rect 11621 15113 11655 15147
rect 12357 15113 12391 15147
rect 12817 15113 12851 15147
rect 16129 15045 16163 15079
rect 3709 14977 3743 15011
rect 3893 14977 3927 15011
rect 4353 14977 4387 15011
rect 5365 14977 5399 15011
rect 9505 14977 9539 15011
rect 10057 14977 10091 15011
rect 10241 14977 10275 15011
rect 11069 14977 11103 15011
rect 11253 14977 11287 15011
rect 11621 14977 11655 15011
rect 11805 14977 11839 15011
rect 12265 14977 12299 15011
rect 12449 14977 12483 15011
rect 12725 14977 12759 15011
rect 13737 14977 13771 15011
rect 16313 14977 16347 15011
rect 16957 14977 16991 15011
rect 1685 14909 1719 14943
rect 1961 14909 1995 14943
rect 3801 14909 3835 14943
rect 4537 14909 4571 14943
rect 5089 14909 5123 14943
rect 6837 14909 6871 14943
rect 7113 14909 7147 14943
rect 9781 14909 9815 14943
rect 15485 14909 15519 14943
rect 5273 14841 5307 14875
rect 13553 14841 13587 14875
rect 3433 14773 3467 14807
rect 4169 14773 4203 14807
rect 5365 14773 5399 14807
rect 16865 14773 16899 14807
rect 5089 14569 5123 14603
rect 6837 14569 6871 14603
rect 8309 14569 8343 14603
rect 14657 14569 14691 14603
rect 15669 14569 15703 14603
rect 16865 14569 16899 14603
rect 5273 14501 5307 14535
rect 12817 14501 12851 14535
rect 6193 14433 6227 14467
rect 9321 14433 9355 14467
rect 9689 14433 9723 14467
rect 9781 14433 9815 14467
rect 11529 14433 11563 14467
rect 13185 14433 13219 14467
rect 16313 14433 16347 14467
rect 1777 14365 1811 14399
rect 4077 14365 4111 14399
rect 4169 14365 4203 14399
rect 4353 14365 4387 14399
rect 4445 14365 4479 14399
rect 6101 14365 6135 14399
rect 6285 14365 6319 14399
rect 6653 14365 6687 14399
rect 7113 14365 7147 14399
rect 7297 14365 7331 14399
rect 7573 14365 7607 14399
rect 8493 14365 8527 14399
rect 9413 14365 9447 14399
rect 9551 14365 9585 14399
rect 10517 14365 10551 14399
rect 10701 14365 10735 14399
rect 10977 14365 11011 14399
rect 11161 14365 11195 14399
rect 11621 14365 11655 14399
rect 12725 14365 12759 14399
rect 12817 14365 12851 14399
rect 12909 14365 12943 14399
rect 13001 14365 13035 14399
rect 13461 14365 13495 14399
rect 14197 14365 14231 14399
rect 14841 14365 14875 14399
rect 15853 14365 15887 14399
rect 16681 14365 16715 14399
rect 2053 14297 2087 14331
rect 4905 14297 4939 14331
rect 5641 14297 5675 14331
rect 13645 14297 13679 14331
rect 3525 14229 3559 14263
rect 3893 14229 3927 14263
rect 5110 14229 5144 14263
rect 5733 14229 5767 14263
rect 7757 14229 7791 14263
rect 9137 14229 9171 14263
rect 10609 14229 10643 14263
rect 11161 14229 11195 14263
rect 11989 14229 12023 14263
rect 14381 14229 14415 14263
rect 15669 14229 15703 14263
rect 2237 14025 2271 14059
rect 3341 14025 3375 14059
rect 7113 14025 7147 14059
rect 2421 13957 2455 13991
rect 6837 13957 6871 13991
rect 9321 13957 9355 13991
rect 11253 13957 11287 13991
rect 14381 13957 14415 13991
rect 2145 13889 2179 13923
rect 4261 13889 4295 13923
rect 4905 13889 4939 13923
rect 5641 13889 5675 13923
rect 5733 13889 5767 13923
rect 5825 13889 5859 13923
rect 6653 13889 6687 13923
rect 7481 13889 7515 13923
rect 8400 13889 8434 13923
rect 8493 13889 8527 13923
rect 8769 13889 8803 13923
rect 8953 13889 8987 13923
rect 9505 13889 9539 13923
rect 10333 13889 10367 13923
rect 10977 13889 11011 13923
rect 11897 13889 11931 13923
rect 14105 13889 14139 13923
rect 16313 13889 16347 13923
rect 2697 13821 2731 13855
rect 2881 13821 2915 13855
rect 2973 13821 3007 13855
rect 4353 13821 4387 13855
rect 4813 13821 4847 13855
rect 6469 13821 6503 13855
rect 7573 13821 7607 13855
rect 7757 13821 7791 13855
rect 10425 13821 10459 13855
rect 11253 13821 11287 13855
rect 11989 13821 12023 13855
rect 12541 13821 12575 13855
rect 12817 13821 12851 13855
rect 15853 13821 15887 13855
rect 2421 13753 2455 13787
rect 5273 13753 5307 13787
rect 8125 13753 8159 13787
rect 11069 13753 11103 13787
rect 16129 13753 16163 13787
rect 3985 13685 4019 13719
rect 6009 13685 6043 13719
rect 8769 13685 8803 13719
rect 10609 13685 10643 13719
rect 12173 13685 12207 13719
rect 2973 13481 3007 13515
rect 7389 13481 7423 13515
rect 8309 13481 8343 13515
rect 11897 13481 11931 13515
rect 13737 13481 13771 13515
rect 15945 13481 15979 13515
rect 16773 13481 16807 13515
rect 4445 13413 4479 13447
rect 3985 13345 4019 13379
rect 5089 13345 5123 13379
rect 6009 13345 6043 13379
rect 7573 13345 7607 13379
rect 10149 13345 10183 13379
rect 13093 13345 13127 13379
rect 13277 13345 13311 13379
rect 14197 13345 14231 13379
rect 14473 13345 14507 13379
rect 3157 13277 3191 13311
rect 3433 13277 3467 13311
rect 4077 13277 4111 13311
rect 4721 13277 4755 13311
rect 4905 13277 4939 13311
rect 5365 13277 5399 13311
rect 5549 13277 5583 13311
rect 5825 13277 5859 13311
rect 6377 13277 6411 13311
rect 6469 13277 6503 13311
rect 6837 13277 6871 13311
rect 7665 13277 7699 13311
rect 8125 13277 8159 13311
rect 8309 13277 8343 13311
rect 9229 13277 9263 13311
rect 9689 13277 9723 13311
rect 9873 13277 9907 13311
rect 13369 13277 13403 13311
rect 16681 13277 16715 13311
rect 3341 13209 3375 13243
rect 7021 13209 7055 13243
rect 10425 13209 10459 13243
rect 9413 13141 9447 13175
rect 9781 13141 9815 13175
rect 6101 12937 6135 12971
rect 7481 12937 7515 12971
rect 8861 12937 8895 12971
rect 10149 12937 10183 12971
rect 10517 12937 10551 12971
rect 10609 12937 10643 12971
rect 11621 12937 11655 12971
rect 15025 12937 15059 12971
rect 15485 12937 15519 12971
rect 3893 12869 3927 12903
rect 5181 12869 5215 12903
rect 7389 12869 7423 12903
rect 9597 12869 9631 12903
rect 9781 12869 9815 12903
rect 12081 12869 12115 12903
rect 3801 12801 3835 12835
rect 3985 12801 4019 12835
rect 4261 12801 4295 12835
rect 4537 12801 4571 12835
rect 5089 12801 5123 12835
rect 5273 12801 5307 12835
rect 5733 12801 5767 12835
rect 6469 12801 6503 12835
rect 6653 12801 6687 12835
rect 8125 12801 8159 12835
rect 9045 12801 9079 12835
rect 14933 12801 14967 12835
rect 15117 12801 15151 12835
rect 15393 12801 15427 12835
rect 15577 12801 15611 12835
rect 16773 12801 16807 12835
rect 16957 12801 16991 12835
rect 17233 12801 17267 12835
rect 17417 12801 17451 12835
rect 4353 12733 4387 12767
rect 5825 12733 5859 12767
rect 6561 12733 6595 12767
rect 7297 12733 7331 12767
rect 10701 12733 10735 12767
rect 7849 12665 7883 12699
rect 11713 12665 11747 12699
rect 4721 12597 4755 12631
rect 8309 12597 8343 12631
rect 16773 12597 16807 12631
rect 17417 12597 17451 12631
rect 10609 12393 10643 12427
rect 13461 12393 13495 12427
rect 17969 12393 18003 12427
rect 4905 12257 4939 12291
rect 17509 12257 17543 12291
rect 19349 12257 19383 12291
rect 2513 12189 2547 12223
rect 2697 12189 2731 12223
rect 4199 12189 4233 12223
rect 4353 12189 4387 12223
rect 4997 12189 5031 12223
rect 5641 12189 5675 12223
rect 9689 12189 9723 12223
rect 9873 12189 9907 12223
rect 11253 12189 11287 12223
rect 11529 12189 11563 12223
rect 13645 12189 13679 12223
rect 14841 12189 14875 12223
rect 15025 12189 15059 12223
rect 17785 12189 17819 12223
rect 18245 12189 18279 12223
rect 18423 12189 18457 12223
rect 18705 12189 18739 12223
rect 18889 12189 18923 12223
rect 10701 12121 10735 12155
rect 17233 12121 17267 12155
rect 19625 12121 19659 12155
rect 2605 12053 2639 12087
rect 3985 12053 4019 12087
rect 5365 12053 5399 12087
rect 5825 12053 5859 12087
rect 9781 12053 9815 12087
rect 11069 12053 11103 12087
rect 11713 12053 11747 12087
rect 14933 12053 14967 12087
rect 15761 12053 15795 12087
rect 18337 12053 18371 12087
rect 18797 12053 18831 12087
rect 21097 12053 21131 12087
rect 9873 11849 9907 11883
rect 10701 11849 10735 11883
rect 11253 11849 11287 11883
rect 11805 11849 11839 11883
rect 15945 11849 15979 11883
rect 17233 11849 17267 11883
rect 20269 11849 20303 11883
rect 5825 11781 5859 11815
rect 8401 11781 8435 11815
rect 11713 11781 11747 11815
rect 12265 11781 12299 11815
rect 3984 11713 4018 11747
rect 4077 11713 4111 11747
rect 6101 11713 6135 11747
rect 8125 11713 8159 11747
rect 10425 11713 10459 11747
rect 11069 11713 11103 11747
rect 11253 11713 11287 11747
rect 13369 11713 13403 11747
rect 16037 11713 16071 11747
rect 16773 11713 16807 11747
rect 17417 11713 17451 11747
rect 17785 11713 17819 11747
rect 20177 11713 20211 11747
rect 1685 11645 1719 11679
rect 1961 11645 1995 11679
rect 10793 11645 10827 11679
rect 13645 11645 13679 11679
rect 15853 11645 15887 11679
rect 18061 11645 18095 11679
rect 20361 11645 20395 11679
rect 3709 11577 3743 11611
rect 12449 11577 12483 11611
rect 16405 11577 16439 11611
rect 19533 11577 19567 11611
rect 3433 11509 3467 11543
rect 4353 11509 4387 11543
rect 10241 11509 10275 11543
rect 15117 11509 15151 11543
rect 16957 11509 16991 11543
rect 19809 11509 19843 11543
rect 2237 11305 2271 11339
rect 4813 11305 4847 11339
rect 6009 11305 6043 11339
rect 6285 11305 6319 11339
rect 9952 11305 9986 11339
rect 11437 11305 11471 11339
rect 11970 11305 12004 11339
rect 14841 11305 14875 11339
rect 17969 11305 18003 11339
rect 19533 11305 19567 11339
rect 21925 11305 21959 11339
rect 2789 11237 2823 11271
rect 7021 11237 7055 11271
rect 7665 11237 7699 11271
rect 14381 11237 14415 11271
rect 18245 11237 18279 11271
rect 20545 11237 20579 11271
rect 22201 11237 22235 11271
rect 3341 11169 3375 11203
rect 4445 11169 4479 11203
rect 5365 11169 5399 11203
rect 5549 11169 5583 11203
rect 9689 11169 9723 11203
rect 11713 11169 11747 11203
rect 16957 11169 16991 11203
rect 17233 11169 17267 11203
rect 18889 11169 18923 11203
rect 21005 11169 21039 11203
rect 21189 11169 21223 11203
rect 22661 11169 22695 11203
rect 22845 11169 22879 11203
rect 2421 11101 2455 11135
rect 3157 11101 3191 11135
rect 4537 11101 4571 11135
rect 6469 11101 6503 11135
rect 6561 11101 6595 11135
rect 6837 11101 6871 11135
rect 7021 11101 7055 11135
rect 7849 11101 7883 11135
rect 8309 11101 8343 11135
rect 9229 11101 9263 11135
rect 9413 11101 9447 11135
rect 14197 11101 14231 11135
rect 17785 11101 17819 11135
rect 18613 11101 18647 11135
rect 19349 11101 19383 11135
rect 20085 11101 20119 11135
rect 21741 11101 21775 11135
rect 6285 11033 6319 11067
rect 9321 11033 9355 11067
rect 14749 11033 14783 11067
rect 18705 11033 18739 11067
rect 22569 11033 22603 11067
rect 3249 10965 3283 10999
rect 5641 10965 5675 10999
rect 8125 10965 8159 10999
rect 13461 10965 13495 10999
rect 15485 10965 15519 10999
rect 20269 10965 20303 10999
rect 20913 10965 20947 10999
rect 3893 10761 3927 10795
rect 4721 10761 4755 10795
rect 7389 10761 7423 10795
rect 10425 10761 10459 10795
rect 10885 10761 10919 10795
rect 11621 10761 11655 10795
rect 12081 10761 12115 10795
rect 13369 10761 13403 10795
rect 13645 10761 13679 10795
rect 15577 10761 15611 10795
rect 16037 10761 16071 10795
rect 3617 10693 3651 10727
rect 8125 10693 8159 10727
rect 9965 10693 9999 10727
rect 12633 10693 12667 10727
rect 14013 10693 14047 10727
rect 22293 10693 22327 10727
rect 2421 10625 2455 10659
rect 2605 10625 2639 10659
rect 3249 10625 3283 10659
rect 3403 10625 3437 10659
rect 4261 10625 4295 10659
rect 5732 10625 5766 10659
rect 5825 10625 5859 10659
rect 6745 10625 6779 10659
rect 7573 10625 7607 10659
rect 7849 10625 7883 10659
rect 9873 10625 9907 10659
rect 10057 10625 10091 10659
rect 10793 10625 10827 10659
rect 11989 10625 12023 10659
rect 12817 10625 12851 10659
rect 13185 10625 13219 10659
rect 14841 10625 14875 10659
rect 15669 10625 15703 10659
rect 16773 10625 16807 10659
rect 17877 10625 17911 10659
rect 21005 10625 21039 10659
rect 21189 10625 21223 10659
rect 4353 10557 4387 10591
rect 5181 10557 5215 10591
rect 6469 10557 6503 10591
rect 11069 10557 11103 10591
rect 12265 10557 12299 10591
rect 14105 10557 14139 10591
rect 14197 10557 14231 10591
rect 15393 10557 15427 10591
rect 18153 10557 18187 10591
rect 22017 10557 22051 10591
rect 4813 10489 4847 10523
rect 6561 10489 6595 10523
rect 9597 10489 9631 10523
rect 2605 10421 2639 10455
rect 5641 10421 5675 10455
rect 6653 10421 6687 10455
rect 14657 10421 14691 10455
rect 16957 10421 16991 10455
rect 19625 10421 19659 10455
rect 21189 10421 21223 10455
rect 23765 10421 23799 10455
rect 5457 10217 5491 10251
rect 6929 10217 6963 10251
rect 7941 10217 7975 10251
rect 9045 10217 9079 10251
rect 12633 10217 12667 10251
rect 14933 10217 14967 10251
rect 16957 10217 16991 10251
rect 19349 10217 19383 10251
rect 22753 10217 22787 10251
rect 4169 10149 4203 10183
rect 7573 10149 7607 10183
rect 16221 10149 16255 10183
rect 4629 10081 4663 10115
rect 4905 10081 4939 10115
rect 8585 10081 8619 10115
rect 9505 10081 9539 10115
rect 9689 10081 9723 10115
rect 10425 10081 10459 10115
rect 15393 10081 15427 10115
rect 15577 10081 15611 10115
rect 17417 10081 17451 10115
rect 17601 10081 17635 10115
rect 18245 10081 18279 10115
rect 20177 10081 20211 10115
rect 23489 10081 23523 10115
rect 23581 10081 23615 10115
rect 1501 10013 1535 10047
rect 4997 10013 5031 10047
rect 5641 10013 5675 10047
rect 5917 10013 5951 10047
rect 6193 10013 6227 10047
rect 6286 10013 6320 10047
rect 6561 10013 6595 10047
rect 6837 10013 6871 10047
rect 7205 10013 7239 10047
rect 7481 10013 7515 10047
rect 7665 10013 7699 10047
rect 9413 10013 9447 10047
rect 12449 10013 12483 10047
rect 12633 10013 12667 10047
rect 13369 10013 13403 10047
rect 14289 10013 14323 10047
rect 16037 10013 16071 10047
rect 18337 10013 18371 10047
rect 18429 10013 18463 10047
rect 19349 10013 19383 10047
rect 19533 10013 19567 10047
rect 22569 10013 22603 10047
rect 22753 10013 22787 10047
rect 1777 9945 1811 9979
rect 3893 9945 3927 9979
rect 8309 9945 8343 9979
rect 10701 9945 10735 9979
rect 14473 9945 14507 9979
rect 17325 9945 17359 9979
rect 20453 9945 20487 9979
rect 23397 9945 23431 9979
rect 3249 9877 3283 9911
rect 4353 9877 4387 9911
rect 5825 9877 5859 9911
rect 6929 9877 6963 9911
rect 7021 9877 7055 9911
rect 8401 9877 8435 9911
rect 12173 9877 12207 9911
rect 13185 9877 13219 9911
rect 15301 9877 15335 9911
rect 18797 9877 18831 9911
rect 21925 9877 21959 9911
rect 23029 9877 23063 9911
rect 2053 9673 2087 9707
rect 2973 9673 3007 9707
rect 9229 9673 9263 9707
rect 10241 9673 10275 9707
rect 15945 9673 15979 9707
rect 18797 9673 18831 9707
rect 3065 9605 3099 9639
rect 6101 9605 6135 9639
rect 6561 9605 6595 9639
rect 11989 9605 12023 9639
rect 14473 9605 14507 9639
rect 17049 9605 17083 9639
rect 2237 9537 2271 9571
rect 4353 9537 4387 9571
rect 4629 9537 4663 9571
rect 4997 9537 5031 9571
rect 5181 9537 5215 9571
rect 5365 9537 5399 9571
rect 5457 9537 5491 9571
rect 5733 9537 5767 9571
rect 5826 9537 5860 9571
rect 6469 9537 6503 9571
rect 6745 9537 6779 9571
rect 7481 9537 7515 9571
rect 10057 9537 10091 9571
rect 10701 9537 10735 9571
rect 11069 9537 11103 9571
rect 11253 9537 11287 9571
rect 11897 9537 11931 9571
rect 12081 9537 12115 9571
rect 18981 9537 19015 9571
rect 19533 9537 19567 9571
rect 22109 9537 22143 9571
rect 22569 9537 22603 9571
rect 23029 9537 23063 9571
rect 3249 9469 3283 9503
rect 7757 9469 7791 9503
rect 14197 9469 14231 9503
rect 16773 9469 16807 9503
rect 18521 9469 18555 9503
rect 19809 9469 19843 9503
rect 21281 9469 21315 9503
rect 23305 9469 23339 9503
rect 24777 9469 24811 9503
rect 2605 9401 2639 9435
rect 4445 9401 4479 9435
rect 4537 9401 4571 9435
rect 11069 9401 11103 9435
rect 22753 9401 22787 9435
rect 4169 9333 4203 9367
rect 5917 9333 5951 9367
rect 6653 9333 6687 9367
rect 10517 9333 10551 9367
rect 22293 9333 22327 9367
rect 6561 9129 6595 9163
rect 7113 9129 7147 9163
rect 7941 9129 7975 9163
rect 11069 9129 11103 9163
rect 15485 9129 15519 9163
rect 17693 9129 17727 9163
rect 23397 9129 23431 9163
rect 24501 9129 24535 9163
rect 3525 9061 3559 9095
rect 4077 9061 4111 9095
rect 6101 9061 6135 9095
rect 15209 9061 15243 9095
rect 21373 9061 21407 9095
rect 3157 8993 3191 9027
rect 4629 8993 4663 9027
rect 5825 8993 5859 9027
rect 9321 8993 9355 9027
rect 9597 8993 9631 9027
rect 13461 8993 13495 9027
rect 14565 8993 14599 9027
rect 19809 8993 19843 9027
rect 19993 8993 20027 9027
rect 22845 8993 22879 9027
rect 23121 8993 23155 9027
rect 23949 8993 23983 9027
rect 2237 8925 2271 8959
rect 3341 8925 3375 8959
rect 5089 8925 5123 8959
rect 5733 8925 5767 8959
rect 6377 8925 6411 8959
rect 6470 8925 6504 8959
rect 7021 8925 7055 8959
rect 7205 8925 7239 8959
rect 8125 8925 8159 8959
rect 14749 8925 14783 8959
rect 15485 8925 15519 8959
rect 15669 8925 15703 8959
rect 16129 8925 16163 8959
rect 17693 8925 17727 8959
rect 17877 8925 17911 8959
rect 19717 8925 19751 8959
rect 24501 8925 24535 8959
rect 24685 8925 24719 8959
rect 4077 8857 4111 8891
rect 13185 8857 13219 8891
rect 20545 8857 20579 8891
rect 2053 8789 2087 8823
rect 4537 8789 4571 8823
rect 4813 8789 4847 8823
rect 5181 8789 5215 8823
rect 6101 8789 6135 8823
rect 7941 8789 7975 8823
rect 11713 8789 11747 8823
rect 14841 8789 14875 8823
rect 15945 8789 15979 8823
rect 19349 8789 19383 8823
rect 20637 8789 20671 8823
rect 21373 8789 21407 8823
rect 23765 8789 23799 8823
rect 23857 8789 23891 8823
rect 3617 8585 3651 8619
rect 4077 8585 4111 8619
rect 10057 8585 10091 8619
rect 10425 8585 10459 8619
rect 10793 8585 10827 8619
rect 11897 8585 11931 8619
rect 12449 8585 12483 8619
rect 12725 8585 12759 8619
rect 13185 8585 13219 8619
rect 17325 8585 17359 8619
rect 17785 8585 17819 8619
rect 18705 8585 18739 8619
rect 19717 8585 19751 8619
rect 20453 8585 20487 8619
rect 22017 8585 22051 8619
rect 1777 8517 1811 8551
rect 4629 8517 4663 8551
rect 7481 8517 7515 8551
rect 9321 8517 9355 8551
rect 9965 8517 9999 8551
rect 15485 8517 15519 8551
rect 3525 8449 3559 8483
rect 4353 8449 4387 8483
rect 4997 8449 5031 8483
rect 5181 8449 5215 8483
rect 5273 8449 5307 8483
rect 5917 8449 5951 8483
rect 7205 8449 7239 8483
rect 9229 8449 9263 8483
rect 9413 8449 9447 8483
rect 10701 8449 10735 8483
rect 10885 8449 10919 8483
rect 11805 8449 11839 8483
rect 11989 8449 12023 8483
rect 12265 8449 12299 8483
rect 13093 8449 13127 8483
rect 17049 8449 17083 8483
rect 17693 8449 17727 8483
rect 18797 8449 18831 8483
rect 19533 8449 19567 8483
rect 20361 8449 20395 8483
rect 20545 8449 20579 8483
rect 20821 8449 20855 8483
rect 21281 8449 21315 8483
rect 21465 8449 21499 8483
rect 21925 8449 21959 8483
rect 22109 8449 22143 8483
rect 23397 8449 23431 8483
rect 1501 8381 1535 8415
rect 3249 8381 3283 8415
rect 4241 8381 4275 8415
rect 4721 8381 4755 8415
rect 6009 8381 6043 8415
rect 9781 8381 9815 8415
rect 13369 8381 13403 8415
rect 14013 8381 14047 8415
rect 15761 8381 15795 8415
rect 17969 8381 18003 8415
rect 18613 8381 18647 8415
rect 23673 8381 23707 8415
rect 4997 8313 5031 8347
rect 5549 8313 5583 8347
rect 8953 8313 8987 8347
rect 19165 8313 19199 8347
rect 16865 8245 16899 8279
rect 21005 8245 21039 8279
rect 21281 8245 21315 8279
rect 25145 8245 25179 8279
rect 2605 8041 2639 8075
rect 4077 8041 4111 8075
rect 4537 8041 4571 8075
rect 6101 8041 6135 8075
rect 10701 8041 10735 8075
rect 12449 8041 12483 8075
rect 14381 8041 14415 8075
rect 15393 8041 15427 8075
rect 23397 8041 23431 8075
rect 23857 8041 23891 8075
rect 2329 7973 2363 8007
rect 5549 7973 5583 8007
rect 9689 7973 9723 8007
rect 24501 7973 24535 8007
rect 3157 7905 3191 7939
rect 8217 7905 8251 7939
rect 10057 7905 10091 7939
rect 10241 7905 10275 7939
rect 16957 7905 16991 7939
rect 21465 7905 21499 7939
rect 21741 7905 21775 7939
rect 24961 7905 24995 7939
rect 25053 7905 25087 7939
rect 2145 7837 2179 7871
rect 2329 7837 2363 7871
rect 2973 7837 3007 7871
rect 3985 7837 4019 7871
rect 4261 7837 4295 7871
rect 4353 7837 4387 7871
rect 5180 7837 5214 7871
rect 5273 7837 5307 7871
rect 5825 7837 5859 7871
rect 6101 7837 6135 7871
rect 6377 7837 6411 7871
rect 7456 7837 7490 7871
rect 8033 7837 8067 7871
rect 8309 7837 8343 7871
rect 12321 7837 12355 7871
rect 12541 7837 12575 7871
rect 12817 7837 12851 7871
rect 13001 7837 13035 7871
rect 14197 7837 14231 7871
rect 14933 7837 14967 7871
rect 15393 7837 15427 7871
rect 15577 7837 15611 7871
rect 15853 7837 15887 7871
rect 16037 7837 16071 7871
rect 16681 7837 16715 7871
rect 18705 7837 18739 7871
rect 18889 7837 18923 7871
rect 19533 7837 19567 7871
rect 23121 7837 23155 7871
rect 23397 7837 23431 7871
rect 23581 7837 23615 7871
rect 24041 7837 24075 7871
rect 24869 7837 24903 7871
rect 5549 7769 5583 7803
rect 6285 7769 6319 7803
rect 9505 7769 9539 7803
rect 15117 7769 15151 7803
rect 18797 7769 18831 7803
rect 3065 7701 3099 7735
rect 4905 7701 4939 7735
rect 5733 7701 5767 7735
rect 7527 7701 7561 7735
rect 7849 7701 7883 7735
rect 10333 7701 10367 7735
rect 12909 7701 12943 7735
rect 15945 7701 15979 7735
rect 18429 7701 18463 7735
rect 19349 7701 19383 7735
rect 19993 7701 20027 7735
rect 22937 7701 22971 7735
rect 4445 7497 4479 7531
rect 6561 7497 6595 7531
rect 7113 7497 7147 7531
rect 20361 7497 20395 7531
rect 20729 7497 20763 7531
rect 21097 7497 21131 7531
rect 21189 7497 21223 7531
rect 24133 7497 24167 7531
rect 3801 7429 3835 7463
rect 8033 7429 8067 7463
rect 16773 7429 16807 7463
rect 18889 7429 18923 7463
rect 22661 7429 22695 7463
rect 2513 7361 2547 7395
rect 2697 7361 2731 7395
rect 4076 7361 4110 7395
rect 4169 7361 4203 7395
rect 4787 7361 4821 7395
rect 5457 7361 5491 7395
rect 6469 7361 6503 7395
rect 6653 7361 6687 7395
rect 7021 7361 7055 7395
rect 7297 7361 7331 7395
rect 9781 7361 9815 7395
rect 11805 7361 11839 7395
rect 12081 7361 12115 7395
rect 12265 7361 12299 7395
rect 15485 7361 15519 7395
rect 16957 7361 16991 7395
rect 19165 7361 19199 7395
rect 19717 7361 19751 7395
rect 19901 7361 19935 7395
rect 20269 7361 20303 7395
rect 20453 7361 20487 7395
rect 21925 7361 21959 7395
rect 22109 7361 22143 7395
rect 22385 7361 22419 7395
rect 24593 7361 24627 7395
rect 4905 7293 4939 7327
rect 5365 7293 5399 7327
rect 7757 7293 7791 7327
rect 13185 7293 13219 7327
rect 13461 7293 13495 7327
rect 15209 7293 15243 7327
rect 17417 7293 17451 7327
rect 21373 7293 21407 7327
rect 5825 7225 5859 7259
rect 24409 7225 24443 7259
rect 2697 7157 2731 7191
rect 7481 7157 7515 7191
rect 9505 7157 9539 7191
rect 9965 7157 9999 7191
rect 11621 7157 11655 7191
rect 12081 7157 12115 7191
rect 14933 7157 14967 7191
rect 21925 7157 21959 7191
rect 3249 6953 3283 6987
rect 6009 6953 6043 6987
rect 8493 6953 8527 6987
rect 9229 6953 9263 6987
rect 11240 6953 11274 6987
rect 13645 6953 13679 6987
rect 18521 6953 18555 6987
rect 23213 6953 23247 6987
rect 24501 6953 24535 6987
rect 1501 6817 1535 6851
rect 5457 6817 5491 6851
rect 7389 6817 7423 6851
rect 9781 6817 9815 6851
rect 10977 6817 11011 6851
rect 15025 6817 15059 6851
rect 20637 6817 20671 6851
rect 23765 6817 23799 6851
rect 25053 6817 25087 6851
rect 4445 6749 4479 6783
rect 4721 6749 4755 6783
rect 5365 6749 5399 6783
rect 5825 6749 5859 6783
rect 6101 6749 6135 6783
rect 7665 6749 7699 6783
rect 7757 6749 7791 6783
rect 7849 6749 7883 6783
rect 8033 6749 8067 6783
rect 9689 6749 9723 6783
rect 9873 6749 9907 6783
rect 13001 6749 13035 6783
rect 13829 6749 13863 6783
rect 14841 6749 14875 6783
rect 15669 6749 15703 6783
rect 17877 6749 17911 6783
rect 18061 6749 18095 6783
rect 18337 6749 18371 6783
rect 20361 6749 20395 6783
rect 23581 6749 23615 6783
rect 24869 6749 24903 6783
rect 1777 6681 1811 6715
rect 4629 6681 4663 6715
rect 5917 6681 5951 6715
rect 8677 6681 8711 6715
rect 9197 6681 9231 6715
rect 9413 6681 9447 6715
rect 3249 6613 3283 6647
rect 4721 6613 4755 6647
rect 4997 6613 5031 6647
rect 8309 6613 8343 6647
rect 8477 6613 8511 6647
rect 9045 6613 9079 6647
rect 12725 6613 12759 6647
rect 13185 6613 13219 6647
rect 14473 6613 14507 6647
rect 14933 6613 14967 6647
rect 15485 6613 15519 6647
rect 17969 6613 18003 6647
rect 22109 6613 22143 6647
rect 23673 6613 23707 6647
rect 24961 6613 24995 6647
rect 2145 6409 2179 6443
rect 2789 6409 2823 6443
rect 3157 6409 3191 6443
rect 6469 6409 6503 6443
rect 8125 6409 8159 6443
rect 9597 6409 9631 6443
rect 11897 6409 11931 6443
rect 12265 6409 12299 6443
rect 20361 6409 20395 6443
rect 20729 6409 20763 6443
rect 21373 6409 21407 6443
rect 21925 6409 21959 6443
rect 25053 6409 25087 6443
rect 7757 6341 7791 6375
rect 13369 6341 13403 6375
rect 18797 6341 18831 6375
rect 7987 6307 8021 6341
rect 2329 6273 2363 6307
rect 4721 6273 4755 6307
rect 5181 6273 5215 6307
rect 5273 6273 5307 6307
rect 5457 6273 5491 6307
rect 5917 6273 5951 6307
rect 6101 6273 6135 6307
rect 6745 6273 6779 6307
rect 8769 6273 8803 6307
rect 9413 6273 9447 6307
rect 9689 6273 9723 6307
rect 9965 6273 9999 6307
rect 10149 6273 10183 6307
rect 11069 6273 11103 6307
rect 13553 6273 13587 6307
rect 16773 6273 16807 6307
rect 17693 6273 17727 6307
rect 17969 6273 18003 6307
rect 18153 6273 18187 6307
rect 18613 6273 18647 6307
rect 20085 6273 20119 6307
rect 21557 6273 21591 6307
rect 22293 6273 22327 6307
rect 23305 6273 23339 6307
rect 3249 6205 3283 6239
rect 3433 6205 3467 6239
rect 4813 6205 4847 6239
rect 5641 6205 5675 6239
rect 6469 6205 6503 6239
rect 8677 6205 8711 6239
rect 12357 6205 12391 6239
rect 12541 6205 12575 6239
rect 14473 6205 14507 6239
rect 14749 6205 14783 6239
rect 20821 6205 20855 6239
rect 20913 6205 20947 6239
rect 22385 6205 22419 6239
rect 22569 6205 22603 6239
rect 23581 6205 23615 6239
rect 4353 6137 4387 6171
rect 6009 6137 6043 6171
rect 6653 6137 6687 6171
rect 10885 6137 10919 6171
rect 7941 6069 7975 6103
rect 8401 6069 8435 6103
rect 9229 6069 9263 6103
rect 10149 6069 10183 6103
rect 16221 6069 16255 6103
rect 16957 6069 16991 6103
rect 17509 6069 17543 6103
rect 18153 6069 18187 6103
rect 18705 6069 18739 6103
rect 19901 6069 19935 6103
rect 5365 5865 5399 5899
rect 7113 5865 7147 5899
rect 11529 5865 11563 5899
rect 15117 5865 15151 5899
rect 23673 5865 23707 5899
rect 2789 5797 2823 5831
rect 6285 5797 6319 5831
rect 7665 5797 7699 5831
rect 13553 5797 13587 5831
rect 15577 5797 15611 5831
rect 4537 5729 4571 5763
rect 4629 5729 4663 5763
rect 5825 5729 5859 5763
rect 12909 5729 12943 5763
rect 16129 5729 16163 5763
rect 19533 5729 19567 5763
rect 19809 5729 19843 5763
rect 2237 5661 2271 5695
rect 2605 5661 2639 5695
rect 2789 5661 2823 5695
rect 3371 5661 3405 5695
rect 3518 5661 3552 5695
rect 4721 5661 4755 5695
rect 4813 5661 4847 5695
rect 5273 5661 5307 5695
rect 5457 5661 5491 5695
rect 5917 5661 5951 5695
rect 6561 5661 6595 5695
rect 6837 5661 6871 5695
rect 7389 5661 7423 5695
rect 7665 5661 7699 5695
rect 7941 5661 7975 5695
rect 8217 5661 8251 5695
rect 8493 5661 8527 5695
rect 9045 5661 9079 5695
rect 11345 5661 11379 5695
rect 12725 5661 12759 5695
rect 15301 5661 15335 5695
rect 16957 5661 16991 5695
rect 23397 5661 23431 5695
rect 23673 5661 23707 5695
rect 23857 5661 23891 5695
rect 6653 5593 6687 5627
rect 7113 5593 7147 5627
rect 8309 5593 8343 5627
rect 8677 5593 8711 5627
rect 9321 5593 9355 5627
rect 12633 5593 12667 5627
rect 13369 5593 13403 5627
rect 17233 5593 17267 5627
rect 2053 5525 2087 5559
rect 3157 5525 3191 5559
rect 4997 5525 5031 5559
rect 6745 5525 6779 5559
rect 7297 5525 7331 5559
rect 7849 5525 7883 5559
rect 10793 5525 10827 5559
rect 11529 5525 11563 5559
rect 12265 5525 12299 5559
rect 15945 5525 15979 5559
rect 16037 5525 16071 5559
rect 18705 5525 18739 5559
rect 21281 5525 21315 5559
rect 23213 5525 23247 5559
rect 3525 5321 3559 5355
rect 3893 5321 3927 5355
rect 3985 5321 4019 5355
rect 6469 5321 6503 5355
rect 7481 5321 7515 5355
rect 8125 5321 8159 5355
rect 10241 5321 10275 5355
rect 15209 5321 15243 5355
rect 15761 5321 15795 5355
rect 16957 5321 16991 5355
rect 17877 5321 17911 5355
rect 18245 5321 18279 5355
rect 18337 5321 18371 5355
rect 20453 5321 20487 5355
rect 21925 5321 21959 5355
rect 22293 5321 22327 5355
rect 1777 5253 1811 5287
rect 4813 5253 4847 5287
rect 5733 5253 5767 5287
rect 7297 5253 7331 5287
rect 9597 5253 9631 5287
rect 13829 5253 13863 5287
rect 1501 5185 1535 5219
rect 4537 5185 4571 5219
rect 4685 5185 4719 5219
rect 4905 5185 4939 5219
rect 5021 5185 5055 5219
rect 6008 5185 6042 5219
rect 6101 5185 6135 5219
rect 6837 5185 6871 5219
rect 7573 5185 7607 5219
rect 10149 5185 10183 5219
rect 10333 5185 10367 5219
rect 11621 5185 11655 5219
rect 14289 5185 14323 5219
rect 14473 5185 14507 5219
rect 15117 5185 15151 5219
rect 16036 5185 16070 5219
rect 16129 5185 16163 5219
rect 16773 5185 16807 5219
rect 19165 5185 19199 5219
rect 20361 5185 20395 5219
rect 20545 5185 20579 5219
rect 21373 5185 21407 5219
rect 23121 5185 23155 5219
rect 3249 5117 3283 5151
rect 4077 5117 4111 5151
rect 6745 5117 6779 5151
rect 9873 5117 9907 5151
rect 11897 5117 11931 5151
rect 15393 5117 15427 5151
rect 18521 5117 18555 5151
rect 19441 5117 19475 5151
rect 22385 5117 22419 5151
rect 22569 5117 22603 5151
rect 23397 5117 23431 5151
rect 5181 5049 5215 5083
rect 7297 5049 7331 5083
rect 14749 5049 14783 5083
rect 16957 5049 16991 5083
rect 8125 4981 8159 5015
rect 13369 4981 13403 5015
rect 13737 4981 13771 5015
rect 14473 4981 14507 5015
rect 21189 4981 21223 5015
rect 24869 4981 24903 5015
rect 2513 4777 2547 4811
rect 2697 4777 2731 4811
rect 4123 4777 4157 4811
rect 7849 4777 7883 4811
rect 8401 4777 8435 4811
rect 9229 4777 9263 4811
rect 11897 4777 11931 4811
rect 12357 4777 12391 4811
rect 16681 4777 16715 4811
rect 22201 4777 22235 4811
rect 23121 4777 23155 4811
rect 23397 4777 23431 4811
rect 4997 4709 5031 4743
rect 5641 4709 5675 4743
rect 6561 4709 6595 4743
rect 10517 4709 10551 4743
rect 16497 4709 16531 4743
rect 24501 4709 24535 4743
rect 2053 4641 2087 4675
rect 3249 4641 3283 4675
rect 4721 4641 4755 4675
rect 6285 4641 6319 4675
rect 7113 4641 7147 4675
rect 14197 4641 14231 4675
rect 19901 4641 19935 4675
rect 20729 4641 20763 4675
rect 23857 4641 23891 4675
rect 24041 4641 24075 4675
rect 24961 4641 24995 4675
rect 25053 4641 25087 4675
rect 1869 4573 1903 4607
rect 3341 4573 3375 4607
rect 4020 4574 4054 4608
rect 4629 4573 4663 4607
rect 5273 4573 5307 4607
rect 5366 4573 5400 4607
rect 6193 4573 6227 4607
rect 7021 4573 7055 4607
rect 7879 4573 7913 4607
rect 8033 4573 8067 4607
rect 8309 4573 8343 4607
rect 8493 4573 8527 4607
rect 9229 4573 9263 4607
rect 9413 4573 9447 4607
rect 12081 4573 12115 4607
rect 12357 4573 12391 4607
rect 12541 4573 12575 4607
rect 12817 4573 12851 4607
rect 13001 4573 13035 4607
rect 13737 4573 13771 4607
rect 17693 4573 17727 4607
rect 18705 4573 18739 4607
rect 19717 4573 19751 4607
rect 20453 4573 20487 4607
rect 22477 4573 22511 4607
rect 22661 4573 22695 4607
rect 22937 4573 22971 4607
rect 2329 4505 2363 4539
rect 2545 4505 2579 4539
rect 10701 4505 10735 4539
rect 13553 4505 13587 4539
rect 14473 4505 14507 4539
rect 16221 4505 16255 4539
rect 2973 4437 3007 4471
rect 7389 4437 7423 4471
rect 12909 4437 12943 4471
rect 15945 4437 15979 4471
rect 17509 4437 17543 4471
rect 18521 4437 18555 4471
rect 19349 4437 19383 4471
rect 19809 4437 19843 4471
rect 22569 4437 22603 4471
rect 23765 4437 23799 4471
rect 24869 4437 24903 4471
rect 4077 4233 4111 4267
rect 4261 4233 4295 4267
rect 6837 4233 6871 4267
rect 10149 4233 10183 4267
rect 17509 4233 17543 4267
rect 17877 4233 17911 4267
rect 24777 4233 24811 4267
rect 8033 4165 8067 4199
rect 18429 4165 18463 4199
rect 1685 4097 1719 4131
rect 3709 4097 3743 4131
rect 4537 4097 4571 4131
rect 4812 4097 4846 4131
rect 4905 4097 4939 4131
rect 7481 4097 7515 4131
rect 7573 4097 7607 4131
rect 7757 4097 7791 4131
rect 8217 4097 8251 4131
rect 8309 4097 8343 4131
rect 9137 4097 9171 4131
rect 9965 4097 9999 4131
rect 10241 4097 10275 4131
rect 10517 4097 10551 4131
rect 10701 4097 10735 4131
rect 10977 4097 11011 4131
rect 11161 4097 11195 4131
rect 11713 4097 11747 4131
rect 14197 4097 14231 4131
rect 14657 4097 14691 4131
rect 20177 4097 20211 4131
rect 20361 4097 20395 4131
rect 20821 4097 20855 4131
rect 21005 4097 21039 4131
rect 23029 4097 23063 4131
rect 1961 4029 1995 4063
rect 3433 4029 3467 4063
rect 6929 4029 6963 4063
rect 7113 4029 7147 4063
rect 9229 4029 9263 4063
rect 9505 4029 9539 4063
rect 11989 4029 12023 4063
rect 14933 4029 14967 4063
rect 17233 4029 17267 4063
rect 17417 4029 17451 4063
rect 18153 4029 18187 4063
rect 20269 4029 20303 4063
rect 23305 4029 23339 4063
rect 14381 3961 14415 3995
rect 16405 3961 16439 3995
rect 21005 3961 21039 3995
rect 4077 3893 4111 3927
rect 6469 3893 6503 3927
rect 7481 3893 7515 3927
rect 8033 3893 8067 3927
rect 9781 3893 9815 3927
rect 10701 3893 10735 3927
rect 11161 3893 11195 3927
rect 13461 3893 13495 3927
rect 19901 3893 19935 3927
rect 2237 3689 2271 3723
rect 2789 3689 2823 3723
rect 6653 3689 6687 3723
rect 7389 3689 7423 3723
rect 10977 3689 11011 3723
rect 12265 3689 12299 3723
rect 16497 3689 16531 3723
rect 18981 3689 19015 3723
rect 23581 3689 23615 3723
rect 12725 3621 12759 3655
rect 20729 3621 20763 3655
rect 5917 3553 5951 3587
rect 7021 3553 7055 3587
rect 9229 3553 9263 3587
rect 13277 3553 13311 3587
rect 17233 3553 17267 3587
rect 17509 3553 17543 3587
rect 21005 3553 21039 3587
rect 22753 3553 22787 3587
rect 2421 3485 2455 3519
rect 2789 3485 2823 3519
rect 2973 3485 3007 3519
rect 4445 3485 4479 3519
rect 4629 3485 4663 3519
rect 6192 3485 6226 3519
rect 6285 3485 6319 3519
rect 6903 3485 6937 3519
rect 7573 3485 7607 3519
rect 7757 3485 7791 3519
rect 7849 3485 7883 3519
rect 8309 3485 8343 3519
rect 8401 3485 8435 3519
rect 8493 3485 8527 3519
rect 12449 3485 12483 3519
rect 13093 3485 13127 3519
rect 14197 3485 14231 3519
rect 16497 3485 16531 3519
rect 16681 3485 16715 3519
rect 19349 3485 19383 3519
rect 19533 3485 19567 3519
rect 20545 3485 20579 3519
rect 20729 3485 20763 3519
rect 23581 3485 23615 3519
rect 23765 3485 23799 3519
rect 9505 3417 9539 3451
rect 19441 3417 19475 3451
rect 22477 3417 22511 3451
rect 4537 3349 4571 3383
rect 8677 3349 8711 3383
rect 13185 3349 13219 3383
rect 14381 3349 14415 3383
rect 3893 3145 3927 3179
rect 5273 3145 5307 3179
rect 7665 3145 7699 3179
rect 8401 3145 8435 3179
rect 11989 3145 12023 3179
rect 15025 3145 15059 3179
rect 15117 3145 15151 3179
rect 17233 3145 17267 3179
rect 21557 3145 21591 3179
rect 22017 3145 22051 3179
rect 4261 3077 4295 3111
rect 4905 3077 4939 3111
rect 5549 3077 5583 3111
rect 9321 3077 9355 3111
rect 17325 3077 17359 3111
rect 3433 3009 3467 3043
rect 3617 3009 3651 3043
rect 4077 3009 4111 3043
rect 4353 3009 4387 3043
rect 5824 3009 5858 3043
rect 5917 3009 5951 3043
rect 6653 3009 6687 3043
rect 7481 3009 7515 3043
rect 7757 3009 7791 3043
rect 8033 3009 8067 3043
rect 8126 3009 8160 3043
rect 9045 3009 9079 3043
rect 12081 3009 12115 3043
rect 12633 3009 12667 3043
rect 12817 3009 12851 3043
rect 13737 3009 13771 3043
rect 14197 3009 14231 3043
rect 14381 3009 14415 3043
rect 16221 3009 16255 3043
rect 16405 3009 16439 3043
rect 19809 3009 19843 3043
rect 21925 3009 21959 3043
rect 22109 3009 22143 3043
rect 4629 2941 4663 2975
rect 4997 2941 5031 2975
rect 5114 2941 5148 2975
rect 6745 2941 6779 2975
rect 12173 2941 12207 2975
rect 15209 2941 15243 2975
rect 17141 2941 17175 2975
rect 20085 2941 20119 2975
rect 3617 2873 3651 2907
rect 7021 2873 7055 2907
rect 13921 2873 13955 2907
rect 7297 2805 7331 2839
rect 10793 2805 10827 2839
rect 11621 2805 11655 2839
rect 12817 2805 12851 2839
rect 14381 2805 14415 2839
rect 14657 2805 14691 2839
rect 16221 2805 16255 2839
rect 17693 2805 17727 2839
rect 8493 2601 8527 2635
rect 14197 2601 14231 2635
rect 16221 2601 16255 2635
rect 3893 2465 3927 2499
rect 5641 2465 5675 2499
rect 7021 2465 7055 2499
rect 7665 2465 7699 2499
rect 10885 2465 10919 2499
rect 15669 2465 15703 2499
rect 15945 2465 15979 2499
rect 19809 2465 19843 2499
rect 19993 2465 20027 2499
rect 3525 2397 3559 2431
rect 5917 2397 5951 2431
rect 6101 2397 6135 2431
rect 7757 2397 7791 2431
rect 8401 2397 8435 2431
rect 8585 2397 8619 2431
rect 13185 2397 13219 2431
rect 13369 2397 13403 2431
rect 13645 2397 13679 2431
rect 13829 2397 13863 2431
rect 17969 2397 18003 2431
rect 18429 2397 18463 2431
rect 18797 2397 18831 2431
rect 20361 2397 20395 2431
rect 20545 2397 20579 2431
rect 4169 2329 4203 2363
rect 6745 2329 6779 2363
rect 11161 2329 11195 2363
rect 13277 2329 13311 2363
rect 17693 2329 17727 2363
rect 3341 2261 3375 2295
rect 6009 2261 6043 2295
rect 6377 2261 6411 2295
rect 6837 2261 6871 2295
rect 8125 2261 8159 2295
rect 12633 2261 12667 2295
rect 13737 2261 13771 2295
rect 18245 2261 18279 2295
rect 18981 2261 19015 2295
rect 19349 2261 19383 2295
rect 19717 2261 19751 2295
rect 20453 2261 20487 2295
rect 4905 2057 4939 2091
rect 5641 2057 5675 2091
rect 7205 2057 7239 2091
rect 9505 2057 9539 2091
rect 12265 2057 12299 2091
rect 12357 2057 12391 2091
rect 13553 2057 13587 2091
rect 18521 2057 18555 2091
rect 3157 1989 3191 2023
rect 6469 1989 6503 2023
rect 13001 1989 13035 2023
rect 15025 1989 15059 2023
rect 19073 1989 19107 2023
rect 2881 1921 2915 1955
rect 5916 1921 5950 1955
rect 6009 1921 6043 1955
rect 6653 1921 6687 1955
rect 7573 1921 7607 1955
rect 8677 1921 8711 1955
rect 11253 1921 11287 1955
rect 12909 1921 12943 1955
rect 13093 1921 13127 1955
rect 15301 1921 15335 1955
rect 16773 1921 16807 1955
rect 4629 1853 4663 1887
rect 5365 1853 5399 1887
rect 6837 1853 6871 1887
rect 6929 1853 6963 1887
rect 7389 1853 7423 1887
rect 7481 1853 7515 1887
rect 7665 1853 7699 1887
rect 8769 1853 8803 1887
rect 10977 1853 11011 1887
rect 12449 1853 12483 1887
rect 17049 1853 17083 1887
rect 18797 1853 18831 1887
rect 5089 1785 5123 1819
rect 8309 1785 8343 1819
rect 11897 1717 11931 1751
rect 13553 1717 13587 1751
rect 20545 1717 20579 1751
rect 4813 1513 4847 1547
rect 6837 1513 6871 1547
rect 8401 1513 8435 1547
rect 11069 1513 11103 1547
rect 11621 1513 11655 1547
rect 17049 1513 17083 1547
rect 9229 1445 9263 1479
rect 1501 1377 1535 1411
rect 7205 1377 7239 1411
rect 7573 1377 7607 1411
rect 8033 1377 8067 1411
rect 15117 1377 15151 1411
rect 18153 1377 18187 1411
rect 3249 1309 3283 1343
rect 4904 1309 4938 1343
rect 4997 1309 5031 1343
rect 7113 1309 7147 1343
rect 7941 1309 7975 1343
rect 8401 1309 8435 1343
rect 8585 1309 8619 1343
rect 9505 1309 9539 1343
rect 11253 1309 11287 1343
rect 11805 1309 11839 1343
rect 14933 1309 14967 1343
rect 17233 1309 17267 1343
rect 17969 1309 18003 1343
rect 15025 1241 15059 1275
rect 18061 1241 18095 1275
rect 9045 1173 9079 1207
rect 14565 1173 14599 1207
rect 17601 1173 17635 1207
<< metal1 >>
rect 1394 21292 1400 21344
rect 1452 21332 1458 21344
rect 13170 21332 13176 21344
rect 1452 21304 13176 21332
rect 1452 21292 1458 21304
rect 13170 21292 13176 21304
rect 13228 21292 13234 21344
rect 3602 21224 3608 21276
rect 3660 21264 3666 21276
rect 14550 21264 14556 21276
rect 3660 21236 14556 21264
rect 3660 21224 3666 21236
rect 14550 21224 14556 21236
rect 14608 21224 14614 21276
rect 5350 21156 5356 21208
rect 5408 21196 5414 21208
rect 14274 21196 14280 21208
rect 5408 21168 14280 21196
rect 5408 21156 5414 21168
rect 14274 21156 14280 21168
rect 14332 21156 14338 21208
rect 9122 20952 9128 21004
rect 9180 20992 9186 21004
rect 9950 20992 9956 21004
rect 9180 20964 9956 20992
rect 9180 20952 9186 20964
rect 9950 20952 9956 20964
rect 10008 20992 10014 21004
rect 15562 20992 15568 21004
rect 10008 20964 15568 20992
rect 10008 20952 10014 20964
rect 15562 20952 15568 20964
rect 15620 20952 15626 21004
rect 7374 20884 7380 20936
rect 7432 20924 7438 20936
rect 15286 20924 15292 20936
rect 7432 20896 15292 20924
rect 7432 20884 7438 20896
rect 15286 20884 15292 20896
rect 15344 20884 15350 20936
rect 9398 20816 9404 20868
rect 9456 20856 9462 20868
rect 14642 20856 14648 20868
rect 9456 20828 14648 20856
rect 9456 20816 9462 20828
rect 14642 20816 14648 20828
rect 14700 20816 14706 20868
rect 11422 20748 11428 20800
rect 11480 20788 11486 20800
rect 14090 20788 14096 20800
rect 11480 20760 14096 20788
rect 11480 20748 11486 20760
rect 14090 20748 14096 20760
rect 14148 20748 14154 20800
rect 1104 20698 25852 20720
rect 1104 20646 8214 20698
rect 8266 20646 8278 20698
rect 8330 20646 8342 20698
rect 8394 20646 8406 20698
rect 8458 20646 8470 20698
rect 8522 20646 16214 20698
rect 16266 20646 16278 20698
rect 16330 20646 16342 20698
rect 16394 20646 16406 20698
rect 16458 20646 16470 20698
rect 16522 20646 24214 20698
rect 24266 20646 24278 20698
rect 24330 20646 24342 20698
rect 24394 20646 24406 20698
rect 24458 20646 24470 20698
rect 24522 20646 25852 20698
rect 1104 20624 25852 20646
rect 5537 20587 5595 20593
rect 5537 20553 5549 20587
rect 5583 20584 5595 20587
rect 8665 20587 8723 20593
rect 5583 20556 6132 20584
rect 5583 20553 5595 20556
rect 5537 20547 5595 20553
rect 4433 20451 4491 20457
rect 4433 20417 4445 20451
rect 4479 20448 4491 20451
rect 4706 20448 4712 20460
rect 4479 20420 4712 20448
rect 4479 20417 4491 20420
rect 4433 20411 4491 20417
rect 4706 20408 4712 20420
rect 4764 20408 4770 20460
rect 4890 20408 4896 20460
rect 4948 20448 4954 20460
rect 5537 20451 5595 20457
rect 5537 20448 5549 20451
rect 4948 20420 5549 20448
rect 4948 20408 4954 20420
rect 5537 20417 5549 20420
rect 5583 20448 5595 20451
rect 5997 20451 6055 20457
rect 5997 20448 6009 20451
rect 5583 20420 6009 20448
rect 5583 20417 5595 20420
rect 5537 20411 5595 20417
rect 5997 20417 6009 20420
rect 6043 20417 6055 20451
rect 6104 20448 6132 20556
rect 8665 20553 8677 20587
rect 8711 20553 8723 20587
rect 8665 20547 8723 20553
rect 8680 20516 8708 20547
rect 8754 20544 8760 20596
rect 8812 20584 8818 20596
rect 10091 20587 10149 20593
rect 10091 20584 10103 20587
rect 8812 20556 10103 20584
rect 8812 20544 8818 20556
rect 10091 20553 10103 20556
rect 10137 20553 10149 20587
rect 10091 20547 10149 20553
rect 12069 20587 12127 20593
rect 12069 20553 12081 20587
rect 12115 20584 12127 20587
rect 14185 20587 14243 20593
rect 12115 20556 12848 20584
rect 12115 20553 12127 20556
rect 12069 20547 12127 20553
rect 9858 20516 9864 20528
rect 8680 20488 9864 20516
rect 9858 20476 9864 20488
rect 9916 20516 9922 20528
rect 9916 20488 10180 20516
rect 9916 20476 9922 20488
rect 6574 20451 6632 20457
rect 6574 20448 6586 20451
rect 6104 20420 6586 20448
rect 5997 20411 6055 20417
rect 6574 20417 6586 20420
rect 6620 20417 6632 20451
rect 6574 20411 6632 20417
rect 7374 20408 7380 20460
rect 7432 20408 7438 20460
rect 7929 20451 7987 20457
rect 7929 20417 7941 20451
rect 7975 20448 7987 20451
rect 8570 20448 8576 20460
rect 7975 20420 8576 20448
rect 7975 20417 7987 20420
rect 7929 20411 7987 20417
rect 8570 20408 8576 20420
rect 8628 20408 8634 20460
rect 9122 20408 9128 20460
rect 9180 20408 9186 20460
rect 9306 20408 9312 20460
rect 9364 20448 9370 20460
rect 10152 20457 10180 20488
rect 11974 20476 11980 20528
rect 12032 20516 12038 20528
rect 12713 20519 12771 20525
rect 12713 20516 12725 20519
rect 12032 20488 12725 20516
rect 12032 20476 12038 20488
rect 12713 20485 12725 20488
rect 12759 20485 12771 20519
rect 12713 20479 12771 20485
rect 9702 20451 9760 20457
rect 9702 20448 9714 20451
rect 9364 20420 9714 20448
rect 9364 20408 9370 20420
rect 9702 20417 9714 20420
rect 9748 20417 9760 20451
rect 10152 20451 10220 20457
rect 10152 20420 10174 20451
rect 9702 20411 9760 20417
rect 10162 20417 10174 20420
rect 10208 20417 10220 20451
rect 12820 20448 12848 20556
rect 14185 20553 14197 20587
rect 14231 20584 14243 20587
rect 16117 20587 16175 20593
rect 14231 20556 15378 20584
rect 14231 20553 14243 20556
rect 14185 20547 14243 20553
rect 10162 20411 10220 20417
rect 12728 20420 12848 20448
rect 12728 20392 12756 20420
rect 13722 20408 13728 20460
rect 13780 20448 13786 20460
rect 14829 20451 14887 20457
rect 14829 20448 14841 20451
rect 13780 20420 14841 20448
rect 13780 20408 13786 20420
rect 14829 20417 14841 20420
rect 14875 20417 14887 20451
rect 15350 20448 15378 20556
rect 16117 20553 16129 20587
rect 16163 20584 16175 20587
rect 16298 20584 16304 20596
rect 16163 20556 16304 20584
rect 16163 20553 16175 20556
rect 16117 20547 16175 20553
rect 16298 20544 16304 20556
rect 16356 20544 16362 20596
rect 15470 20457 15476 20460
rect 15422 20452 15476 20457
rect 15421 20451 15476 20452
rect 15421 20448 15434 20451
rect 15350 20420 15434 20448
rect 14829 20411 14887 20417
rect 15422 20417 15434 20420
rect 15468 20417 15476 20451
rect 15422 20411 15476 20417
rect 15470 20408 15476 20411
rect 15528 20408 15534 20460
rect 198 20340 204 20392
rect 256 20380 262 20392
rect 4617 20383 4675 20389
rect 4617 20380 4629 20383
rect 256 20352 4629 20380
rect 256 20340 262 20352
rect 4617 20349 4629 20352
rect 4663 20349 4675 20383
rect 4617 20343 4675 20349
rect 5166 20340 5172 20392
rect 5224 20340 5230 20392
rect 8297 20383 8355 20389
rect 8297 20349 8309 20383
rect 8343 20380 8355 20383
rect 10042 20380 10048 20392
rect 8343 20352 10048 20380
rect 8343 20349 8355 20352
rect 8297 20343 8355 20349
rect 10042 20340 10048 20352
rect 10100 20380 10106 20392
rect 11146 20380 11152 20392
rect 10100 20352 11152 20380
rect 10100 20340 10106 20352
rect 11146 20340 11152 20352
rect 11204 20340 11210 20392
rect 11238 20340 11244 20392
rect 11296 20380 11302 20392
rect 11701 20383 11759 20389
rect 11701 20380 11713 20383
rect 11296 20352 11713 20380
rect 11296 20340 11302 20352
rect 11701 20349 11713 20352
rect 11747 20380 11759 20383
rect 12345 20383 12403 20389
rect 12345 20380 12357 20383
rect 11747 20352 12357 20380
rect 11747 20349 11759 20352
rect 11701 20343 11759 20349
rect 12345 20349 12357 20352
rect 12391 20349 12403 20383
rect 12345 20343 12403 20349
rect 12710 20340 12716 20392
rect 12768 20340 12774 20392
rect 13630 20340 13636 20392
rect 13688 20380 13694 20392
rect 14553 20383 14611 20389
rect 14553 20380 14565 20383
rect 13688 20352 14565 20380
rect 13688 20340 13694 20352
rect 14553 20349 14565 20352
rect 14599 20380 14611 20383
rect 15654 20380 15660 20392
rect 14599 20352 15660 20380
rect 14599 20349 14611 20352
rect 14553 20343 14611 20349
rect 15654 20340 15660 20352
rect 15712 20340 15718 20392
rect 15746 20340 15752 20392
rect 15804 20340 15810 20392
rect 8665 20315 8723 20321
rect 8665 20281 8677 20315
rect 8711 20312 8723 20315
rect 10226 20312 10232 20324
rect 8711 20284 10232 20312
rect 8711 20281 8723 20284
rect 8665 20275 8723 20281
rect 10226 20272 10232 20284
rect 10284 20272 10290 20324
rect 12066 20272 12072 20324
rect 12124 20272 12130 20324
rect 14182 20272 14188 20324
rect 14240 20272 14246 20324
rect 16117 20315 16175 20321
rect 16117 20281 16129 20315
rect 16163 20312 16175 20315
rect 17218 20312 17224 20324
rect 16163 20284 17224 20312
rect 16163 20281 16175 20284
rect 16117 20275 16175 20281
rect 17218 20272 17224 20284
rect 17276 20272 17282 20324
rect 5350 20204 5356 20256
rect 5408 20204 5414 20256
rect 5534 20204 5540 20256
rect 5592 20244 5598 20256
rect 5813 20247 5871 20253
rect 5813 20244 5825 20247
rect 5592 20216 5825 20244
rect 5592 20204 5598 20216
rect 5813 20213 5825 20216
rect 5859 20213 5871 20247
rect 5813 20207 5871 20213
rect 5902 20204 5908 20256
rect 5960 20244 5966 20256
rect 6503 20247 6561 20253
rect 6503 20244 6515 20247
rect 5960 20216 6515 20244
rect 5960 20204 5966 20216
rect 6503 20213 6515 20216
rect 6549 20213 6561 20247
rect 6503 20207 6561 20213
rect 7377 20247 7435 20253
rect 7377 20213 7389 20247
rect 7423 20244 7435 20247
rect 7466 20244 7472 20256
rect 7423 20216 7472 20244
rect 7423 20213 7435 20216
rect 7377 20207 7435 20213
rect 7466 20204 7472 20216
rect 7524 20204 7530 20256
rect 9309 20247 9367 20253
rect 9309 20213 9321 20247
rect 9355 20244 9367 20247
rect 9398 20244 9404 20256
rect 9355 20216 9404 20244
rect 9355 20213 9367 20216
rect 9309 20207 9367 20213
rect 9398 20204 9404 20216
rect 9456 20204 9462 20256
rect 9490 20204 9496 20256
rect 9548 20244 9554 20256
rect 9631 20247 9689 20253
rect 9631 20244 9643 20247
rect 9548 20216 9643 20244
rect 9548 20204 9554 20216
rect 9631 20213 9643 20216
rect 9677 20213 9689 20247
rect 9631 20207 9689 20213
rect 12710 20204 12716 20256
rect 12768 20204 12774 20256
rect 15010 20204 15016 20256
rect 15068 20204 15074 20256
rect 15194 20204 15200 20256
rect 15252 20244 15258 20256
rect 15335 20247 15393 20253
rect 15335 20244 15347 20247
rect 15252 20216 15347 20244
rect 15252 20204 15258 20216
rect 15335 20213 15347 20216
rect 15381 20213 15393 20247
rect 15335 20207 15393 20213
rect 1104 20154 25852 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 12214 20154
rect 12266 20102 12278 20154
rect 12330 20102 12342 20154
rect 12394 20102 12406 20154
rect 12458 20102 12470 20154
rect 12522 20102 20214 20154
rect 20266 20102 20278 20154
rect 20330 20102 20342 20154
rect 20394 20102 20406 20154
rect 20458 20102 20470 20154
rect 20522 20102 25852 20154
rect 1104 20080 25852 20102
rect 6181 20043 6239 20049
rect 6181 20009 6193 20043
rect 6227 20040 6239 20043
rect 6227 20012 9812 20040
rect 6227 20009 6239 20012
rect 6181 20003 6239 20009
rect 4801 19975 4859 19981
rect 4801 19941 4813 19975
rect 4847 19972 4859 19975
rect 5537 19975 5595 19981
rect 5537 19972 5549 19975
rect 4847 19944 5549 19972
rect 4847 19941 4859 19944
rect 4801 19935 4859 19941
rect 5537 19941 5549 19944
rect 5583 19941 5595 19975
rect 5537 19935 5595 19941
rect 7745 19975 7803 19981
rect 7745 19941 7757 19975
rect 7791 19972 7803 19975
rect 8481 19975 8539 19981
rect 8481 19972 8493 19975
rect 7791 19944 8493 19972
rect 7791 19941 7803 19944
rect 7745 19935 7803 19941
rect 8481 19941 8493 19944
rect 8527 19941 8539 19975
rect 8481 19935 8539 19941
rect 9398 19932 9404 19984
rect 9456 19932 9462 19984
rect 9784 19972 9812 20012
rect 9858 20000 9864 20052
rect 9916 20000 9922 20052
rect 11974 20040 11980 20052
rect 9968 20012 11980 20040
rect 9968 19972 9996 20012
rect 11974 20000 11980 20012
rect 12032 20000 12038 20052
rect 12066 20000 12072 20052
rect 12124 20040 12130 20052
rect 12161 20043 12219 20049
rect 12161 20040 12173 20043
rect 12124 20012 12173 20040
rect 12124 20000 12130 20012
rect 12161 20009 12173 20012
rect 12207 20009 12219 20043
rect 13446 20040 13452 20052
rect 12161 20003 12219 20009
rect 12268 20012 13452 20040
rect 9784 19944 9996 19972
rect 10321 19975 10379 19981
rect 10321 19941 10333 19975
rect 10367 19941 10379 19975
rect 10321 19935 10379 19941
rect 5629 19907 5687 19913
rect 5629 19873 5641 19907
rect 5675 19904 5687 19907
rect 5902 19904 5908 19916
rect 5675 19876 5908 19904
rect 5675 19873 5687 19876
rect 5629 19867 5687 19873
rect 5902 19864 5908 19876
rect 5960 19864 5966 19916
rect 7561 19907 7619 19913
rect 7561 19904 7573 19907
rect 6748 19876 7573 19904
rect 4249 19839 4307 19845
rect 4249 19805 4261 19839
rect 4295 19805 4307 19839
rect 4249 19799 4307 19805
rect 4801 19839 4859 19845
rect 4801 19805 4813 19839
rect 4847 19836 4859 19839
rect 4890 19836 4896 19848
rect 4847 19808 4896 19836
rect 4847 19805 4859 19808
rect 4801 19799 4859 19805
rect 4264 19768 4292 19799
rect 4890 19796 4896 19808
rect 4948 19796 4954 19848
rect 5077 19839 5135 19845
rect 5077 19805 5089 19839
rect 5123 19836 5135 19839
rect 5442 19836 5448 19848
rect 5123 19808 5448 19836
rect 5123 19805 5135 19808
rect 5077 19799 5135 19805
rect 5092 19768 5120 19799
rect 5442 19796 5448 19808
rect 5500 19796 5506 19848
rect 6748 19845 6776 19876
rect 7561 19873 7573 19876
rect 7607 19873 7619 19907
rect 8021 19907 8079 19913
rect 8021 19904 8033 19907
rect 7561 19867 7619 19873
rect 7668 19876 8033 19904
rect 5537 19839 5595 19845
rect 5537 19805 5549 19839
rect 5583 19836 5595 19839
rect 5997 19839 6055 19845
rect 5997 19836 6009 19839
rect 5583 19808 6009 19836
rect 5583 19805 5595 19808
rect 5537 19799 5595 19805
rect 5997 19805 6009 19808
rect 6043 19805 6055 19839
rect 5997 19799 6055 19805
rect 6733 19839 6791 19845
rect 6733 19805 6745 19839
rect 6779 19805 6791 19839
rect 6733 19799 6791 19805
rect 7006 19796 7012 19848
rect 7064 19836 7070 19848
rect 7193 19839 7251 19845
rect 7193 19836 7205 19839
rect 7064 19808 7205 19836
rect 7064 19796 7070 19808
rect 7193 19805 7205 19808
rect 7239 19836 7251 19839
rect 7668 19836 7696 19876
rect 8021 19873 8033 19876
rect 8067 19873 8079 19907
rect 8021 19867 8079 19873
rect 8573 19907 8631 19913
rect 8573 19873 8585 19907
rect 8619 19904 8631 19907
rect 9490 19904 9496 19916
rect 8619 19876 9496 19904
rect 8619 19873 8631 19876
rect 8573 19867 8631 19873
rect 9490 19864 9496 19876
rect 9548 19864 9554 19916
rect 10042 19864 10048 19916
rect 10100 19864 10106 19916
rect 10226 19864 10232 19916
rect 10284 19904 10290 19916
rect 10336 19904 10364 19935
rect 11146 19932 11152 19984
rect 11204 19932 11210 19984
rect 12268 19972 12296 20012
rect 13446 20000 13452 20012
rect 13504 20000 13510 20052
rect 14182 20000 14188 20052
rect 14240 20000 14246 20052
rect 15378 20040 15384 20052
rect 14292 20012 15384 20040
rect 11256 19944 12296 19972
rect 12437 19975 12495 19981
rect 10284 19876 10364 19904
rect 10284 19864 10290 19876
rect 10410 19864 10416 19916
rect 10468 19904 10474 19916
rect 11256 19904 11284 19944
rect 12437 19941 12449 19975
rect 12483 19972 12495 19975
rect 13722 19972 13728 19984
rect 12483 19944 13728 19972
rect 12483 19941 12495 19944
rect 12437 19935 12495 19941
rect 13722 19932 13728 19944
rect 13780 19932 13786 19984
rect 14292 19904 14320 20012
rect 15378 20000 15384 20012
rect 15436 20000 15442 20052
rect 15470 20000 15476 20052
rect 15528 20000 15534 20052
rect 16298 20000 16304 20052
rect 16356 20000 16362 20052
rect 17218 20000 17224 20052
rect 17276 20000 17282 20052
rect 15010 19932 15016 19984
rect 15068 19972 15074 19984
rect 16485 19975 16543 19981
rect 15068 19944 15516 19972
rect 15068 19932 15074 19944
rect 15028 19904 15056 19932
rect 10468 19876 11284 19904
rect 11348 19876 14320 19904
rect 14384 19876 15056 19904
rect 10468 19864 10474 19876
rect 7239 19808 7696 19836
rect 7745 19839 7803 19845
rect 7239 19805 7251 19808
rect 7193 19799 7251 19805
rect 7745 19805 7757 19839
rect 7791 19836 7803 19839
rect 8938 19836 8944 19848
rect 7791 19808 8944 19836
rect 7791 19805 7803 19808
rect 7745 19799 7803 19805
rect 8938 19796 8944 19808
rect 8996 19796 9002 19848
rect 9033 19839 9091 19845
rect 9033 19805 9045 19839
rect 9079 19836 9091 19839
rect 9122 19836 9128 19848
rect 9079 19808 9128 19836
rect 9079 19805 9091 19808
rect 9033 19799 9091 19805
rect 9122 19796 9128 19808
rect 9180 19796 9186 19848
rect 11348 19845 11376 19876
rect 9677 19839 9735 19845
rect 9677 19805 9689 19839
rect 9723 19836 9735 19839
rect 10505 19839 10563 19845
rect 10505 19836 10517 19839
rect 9723 19808 10517 19836
rect 9723 19805 9735 19808
rect 9677 19799 9735 19805
rect 10505 19805 10517 19808
rect 10551 19805 10563 19839
rect 10505 19799 10563 19805
rect 11333 19839 11391 19845
rect 11333 19805 11345 19839
rect 11379 19805 11391 19839
rect 11333 19799 11391 19805
rect 7374 19768 7380 19780
rect 4264 19740 5120 19768
rect 6932 19740 7380 19768
rect 6932 19709 6960 19740
rect 7374 19728 7380 19740
rect 7432 19768 7438 19780
rect 9692 19768 9720 19799
rect 11606 19796 11612 19848
rect 11664 19836 11670 19848
rect 11701 19839 11759 19845
rect 11701 19836 11713 19839
rect 11664 19808 11713 19836
rect 11664 19796 11670 19808
rect 11701 19805 11713 19808
rect 11747 19805 11759 19839
rect 11701 19799 11759 19805
rect 11974 19796 11980 19848
rect 12032 19836 12038 19848
rect 12437 19839 12495 19845
rect 12437 19836 12449 19839
rect 12032 19808 12449 19836
rect 12032 19796 12038 19808
rect 12437 19805 12449 19808
rect 12483 19805 12495 19839
rect 12437 19799 12495 19805
rect 12986 19796 12992 19848
rect 13044 19836 13050 19848
rect 14384 19845 14412 19876
rect 15194 19864 15200 19916
rect 15252 19864 15258 19916
rect 15488 19913 15516 19944
rect 16485 19941 16497 19975
rect 16531 19941 16543 19975
rect 16485 19935 16543 19941
rect 15473 19907 15531 19913
rect 15473 19873 15485 19907
rect 15519 19873 15531 19907
rect 15473 19867 15531 19873
rect 15654 19864 15660 19916
rect 15712 19904 15718 19916
rect 15841 19907 15899 19913
rect 15841 19904 15853 19907
rect 15712 19876 15853 19904
rect 15712 19864 15718 19876
rect 15841 19873 15853 19876
rect 15887 19873 15899 19907
rect 15841 19867 15899 19873
rect 13265 19839 13323 19845
rect 13265 19836 13277 19839
rect 13044 19808 13277 19836
rect 13044 19796 13050 19808
rect 13265 19805 13277 19808
rect 13311 19805 13323 19839
rect 13265 19799 13323 19805
rect 14369 19839 14427 19845
rect 14369 19805 14381 19839
rect 14415 19805 14427 19839
rect 14369 19799 14427 19805
rect 14645 19839 14703 19845
rect 14645 19805 14657 19839
rect 14691 19805 14703 19839
rect 14645 19799 14703 19805
rect 16117 19839 16175 19845
rect 16117 19805 16129 19839
rect 16163 19805 16175 19839
rect 16500 19836 16528 19935
rect 16666 19932 16672 19984
rect 16724 19972 16730 19984
rect 24854 19972 24860 19984
rect 16724 19944 24860 19972
rect 16724 19932 16730 19944
rect 24854 19932 24860 19944
rect 24912 19932 24918 19984
rect 16878 19839 16936 19845
rect 16878 19836 16890 19839
rect 16500 19808 16890 19836
rect 16117 19799 16175 19805
rect 16878 19805 16890 19808
rect 16924 19805 16936 19839
rect 16878 19799 16936 19805
rect 17405 19839 17463 19845
rect 17405 19805 17417 19839
rect 17451 19805 17463 19839
rect 17405 19799 17463 19805
rect 7432 19740 9720 19768
rect 7432 19728 7438 19740
rect 11422 19728 11428 19780
rect 11480 19728 11486 19780
rect 11517 19771 11575 19777
rect 11517 19737 11529 19771
rect 11563 19737 11575 19771
rect 11517 19731 11575 19737
rect 6917 19703 6975 19709
rect 6917 19669 6929 19703
rect 6963 19669 6975 19703
rect 6917 19663 6975 19669
rect 9398 19660 9404 19712
rect 9456 19660 9462 19712
rect 10870 19660 10876 19712
rect 10928 19700 10934 19712
rect 11532 19700 11560 19731
rect 13814 19728 13820 19780
rect 13872 19728 13878 19780
rect 14182 19728 14188 19780
rect 14240 19768 14246 19780
rect 14660 19768 14688 19799
rect 14240 19740 14688 19768
rect 15105 19771 15163 19777
rect 14240 19728 14246 19740
rect 15105 19737 15117 19771
rect 15151 19768 15163 19771
rect 15470 19768 15476 19780
rect 15151 19740 15476 19768
rect 15151 19737 15163 19740
rect 15105 19731 15163 19737
rect 15470 19728 15476 19740
rect 15528 19728 15534 19780
rect 10928 19672 11560 19700
rect 10928 19660 10934 19672
rect 12250 19660 12256 19712
rect 12308 19700 12314 19712
rect 15746 19700 15752 19712
rect 12308 19672 15752 19700
rect 12308 19660 12314 19672
rect 15746 19660 15752 19672
rect 15804 19700 15810 19712
rect 16132 19700 16160 19799
rect 16485 19771 16543 19777
rect 16485 19737 16497 19771
rect 16531 19768 16543 19771
rect 16574 19768 16580 19780
rect 16531 19740 16580 19768
rect 16531 19737 16543 19740
rect 16485 19731 16543 19737
rect 16574 19728 16580 19740
rect 16632 19768 16638 19780
rect 17420 19768 17448 19799
rect 16632 19740 17448 19768
rect 16632 19728 16638 19740
rect 15804 19672 16160 19700
rect 15804 19660 15810 19672
rect 16758 19660 16764 19712
rect 16816 19709 16822 19712
rect 16816 19703 16865 19709
rect 16816 19669 16819 19703
rect 16853 19669 16865 19703
rect 16816 19663 16865 19669
rect 16816 19660 16822 19663
rect 1104 19610 25852 19632
rect 1104 19558 8214 19610
rect 8266 19558 8278 19610
rect 8330 19558 8342 19610
rect 8394 19558 8406 19610
rect 8458 19558 8470 19610
rect 8522 19558 16214 19610
rect 16266 19558 16278 19610
rect 16330 19558 16342 19610
rect 16394 19558 16406 19610
rect 16458 19558 16470 19610
rect 16522 19558 24214 19610
rect 24266 19558 24278 19610
rect 24330 19558 24342 19610
rect 24394 19558 24406 19610
rect 24458 19558 24470 19610
rect 24522 19558 25852 19610
rect 1104 19536 25852 19558
rect 5350 19456 5356 19508
rect 5408 19456 5414 19508
rect 5442 19456 5448 19508
rect 5500 19496 5506 19508
rect 5721 19499 5779 19505
rect 5721 19496 5733 19499
rect 5500 19468 5733 19496
rect 5500 19456 5506 19468
rect 5721 19465 5733 19468
rect 5767 19465 5779 19499
rect 5721 19459 5779 19465
rect 7006 19456 7012 19508
rect 7064 19456 7070 19508
rect 9398 19456 9404 19508
rect 9456 19496 9462 19508
rect 9953 19499 10011 19505
rect 9953 19496 9965 19499
rect 9456 19468 9965 19496
rect 9456 19456 9462 19468
rect 9953 19465 9965 19468
rect 9999 19465 10011 19499
rect 9953 19459 10011 19465
rect 11238 19456 11244 19508
rect 11296 19456 11302 19508
rect 12250 19456 12256 19508
rect 12308 19456 12314 19508
rect 13127 19499 13185 19505
rect 13127 19465 13139 19499
rect 13173 19496 13185 19499
rect 13814 19496 13820 19508
rect 13173 19468 13820 19496
rect 13173 19465 13185 19468
rect 13127 19459 13185 19465
rect 13814 19456 13820 19468
rect 13872 19456 13878 19508
rect 16393 19499 16451 19505
rect 14660 19468 15516 19496
rect 4433 19431 4491 19437
rect 4433 19397 4445 19431
rect 4479 19428 4491 19431
rect 4706 19428 4712 19440
rect 4479 19400 4712 19428
rect 4479 19397 4491 19400
rect 4433 19391 4491 19397
rect 4706 19388 4712 19400
rect 4764 19388 4770 19440
rect 7745 19431 7803 19437
rect 7745 19397 7757 19431
rect 7791 19428 7803 19431
rect 8754 19428 8760 19440
rect 7791 19400 8760 19428
rect 7791 19397 7803 19400
rect 7745 19391 7803 19397
rect 8754 19388 8760 19400
rect 8812 19388 8818 19440
rect 9217 19431 9275 19437
rect 9217 19397 9229 19431
rect 9263 19428 9275 19431
rect 10042 19428 10048 19440
rect 9263 19400 10048 19428
rect 9263 19397 9275 19400
rect 9217 19391 9275 19397
rect 10042 19388 10048 19400
rect 10100 19388 10106 19440
rect 10778 19437 10784 19440
rect 10755 19431 10784 19437
rect 10755 19397 10767 19431
rect 10755 19391 10784 19397
rect 10778 19388 10784 19391
rect 10836 19388 10842 19440
rect 10965 19431 11023 19437
rect 10965 19397 10977 19431
rect 11011 19428 11023 19431
rect 11606 19428 11612 19440
rect 11011 19400 11612 19428
rect 11011 19397 11023 19400
rect 10965 19391 11023 19397
rect 11606 19388 11612 19400
rect 11664 19388 11670 19440
rect 14660 19437 14688 19468
rect 15488 19440 15516 19468
rect 16393 19465 16405 19499
rect 16439 19496 16451 19499
rect 16574 19496 16580 19508
rect 16439 19468 16580 19496
rect 16439 19465 16451 19468
rect 16393 19459 16451 19465
rect 11767 19431 11825 19437
rect 11767 19397 11779 19431
rect 11813 19428 11825 19431
rect 12529 19431 12587 19437
rect 12529 19428 12541 19431
rect 11813 19400 12541 19428
rect 11813 19397 11825 19400
rect 11767 19391 11825 19397
rect 12529 19397 12541 19400
rect 12575 19397 12587 19431
rect 12529 19391 12587 19397
rect 14645 19431 14703 19437
rect 14645 19397 14657 19431
rect 14691 19397 14703 19431
rect 14645 19391 14703 19397
rect 15381 19385 15439 19391
rect 15470 19388 15476 19440
rect 15528 19428 15534 19440
rect 15528 19400 16252 19428
rect 15528 19388 15534 19400
rect 4341 19363 4399 19369
rect 4341 19329 4353 19363
rect 4387 19360 4399 19363
rect 4798 19360 4804 19372
rect 4387 19332 4804 19360
rect 4387 19329 4399 19332
rect 4341 19323 4399 19329
rect 4798 19320 4804 19332
rect 4856 19320 4862 19372
rect 5810 19320 5816 19372
rect 5868 19320 5874 19372
rect 6825 19363 6883 19369
rect 6825 19329 6837 19363
rect 6871 19360 6883 19363
rect 7098 19360 7104 19372
rect 6871 19332 7104 19360
rect 6871 19329 6883 19332
rect 6825 19323 6883 19329
rect 7098 19320 7104 19332
rect 7156 19320 7162 19372
rect 7466 19320 7472 19372
rect 7524 19360 7530 19372
rect 7837 19363 7895 19369
rect 7837 19360 7849 19363
rect 7524 19332 7849 19360
rect 7524 19320 7530 19332
rect 7837 19329 7849 19332
rect 7883 19329 7895 19363
rect 7837 19323 7895 19329
rect 8297 19363 8355 19369
rect 8297 19329 8309 19363
rect 8343 19360 8355 19363
rect 8570 19360 8576 19372
rect 8343 19332 8576 19360
rect 8343 19329 8355 19332
rect 8297 19323 8355 19329
rect 8570 19320 8576 19332
rect 8628 19320 8634 19372
rect 9030 19320 9036 19372
rect 9088 19320 9094 19372
rect 9309 19363 9367 19369
rect 9309 19329 9321 19363
rect 9355 19360 9367 19363
rect 10410 19360 10416 19372
rect 9355 19332 10416 19360
rect 9355 19329 9367 19332
rect 9309 19323 9367 19329
rect 10410 19320 10416 19332
rect 10468 19320 10474 19372
rect 10870 19320 10876 19372
rect 10928 19320 10934 19372
rect 11054 19320 11060 19372
rect 11112 19320 11118 19372
rect 11514 19320 11520 19372
rect 11572 19360 11578 19372
rect 11885 19363 11943 19369
rect 11885 19360 11897 19363
rect 11572 19332 11897 19360
rect 11572 19320 11578 19332
rect 11885 19329 11897 19332
rect 11931 19329 11943 19363
rect 11885 19323 11943 19329
rect 11977 19363 12035 19369
rect 11977 19329 11989 19363
rect 12023 19329 12035 19363
rect 11977 19323 12035 19329
rect 4985 19295 5043 19301
rect 4985 19261 4997 19295
rect 5031 19261 5043 19295
rect 4985 19255 5043 19261
rect 5353 19295 5411 19301
rect 5353 19261 5365 19295
rect 5399 19292 5411 19295
rect 5534 19292 5540 19304
rect 5399 19264 5540 19292
rect 5399 19261 5411 19264
rect 5353 19255 5411 19261
rect 5000 19224 5028 19255
rect 5534 19252 5540 19264
rect 5592 19252 5598 19304
rect 8849 19295 8907 19301
rect 8849 19261 8861 19295
rect 8895 19292 8907 19295
rect 9122 19292 9128 19304
rect 8895 19264 9128 19292
rect 8895 19261 8907 19264
rect 8849 19255 8907 19261
rect 9122 19252 9128 19264
rect 9180 19292 9186 19304
rect 9585 19295 9643 19301
rect 9585 19292 9597 19295
rect 9180 19264 9597 19292
rect 9180 19252 9186 19264
rect 9585 19261 9597 19264
rect 9631 19261 9643 19295
rect 9585 19255 9643 19261
rect 9950 19252 9956 19304
rect 10008 19252 10014 19304
rect 10597 19295 10655 19301
rect 10597 19261 10609 19295
rect 10643 19292 10655 19295
rect 11238 19292 11244 19304
rect 10643 19264 11244 19292
rect 10643 19261 10655 19264
rect 10597 19255 10655 19261
rect 5166 19224 5172 19236
rect 5000 19196 5172 19224
rect 5166 19184 5172 19196
rect 5224 19224 5230 19236
rect 5224 19196 7420 19224
rect 5224 19184 5230 19196
rect 7282 19116 7288 19168
rect 7340 19116 7346 19168
rect 7392 19156 7420 19196
rect 9490 19184 9496 19236
rect 9548 19224 9554 19236
rect 10612 19224 10640 19255
rect 11238 19252 11244 19264
rect 11296 19292 11302 19304
rect 11422 19292 11428 19304
rect 11296 19264 11428 19292
rect 11296 19252 11302 19264
rect 11422 19252 11428 19264
rect 11480 19292 11486 19304
rect 11609 19295 11667 19301
rect 11609 19292 11621 19295
rect 11480 19264 11621 19292
rect 11480 19252 11486 19264
rect 11609 19261 11621 19264
rect 11655 19261 11667 19295
rect 11609 19255 11667 19261
rect 9548 19196 10640 19224
rect 9548 19184 9554 19196
rect 10870 19184 10876 19236
rect 10928 19224 10934 19236
rect 11992 19224 12020 19323
rect 12066 19320 12072 19372
rect 12124 19320 12130 19372
rect 12710 19320 12716 19372
rect 12768 19360 12774 19372
rect 13024 19363 13082 19369
rect 13024 19360 13036 19363
rect 12768 19332 13036 19360
rect 12768 19320 12774 19332
rect 13024 19329 13036 19332
rect 13070 19329 13082 19363
rect 13024 19323 13082 19329
rect 14182 19320 14188 19372
rect 14240 19320 14246 19372
rect 14737 19363 14795 19369
rect 14737 19329 14749 19363
rect 14783 19360 14795 19363
rect 15010 19360 15016 19372
rect 14783 19332 15016 19360
rect 14783 19329 14795 19332
rect 14737 19323 14795 19329
rect 15010 19320 15016 19332
rect 15068 19320 15074 19372
rect 15381 19351 15393 19385
rect 15427 19351 15439 19385
rect 16224 19369 16252 19400
rect 15381 19345 15439 19351
rect 15933 19363 15991 19369
rect 15396 19304 15424 19345
rect 15933 19329 15945 19363
rect 15979 19360 15991 19363
rect 16209 19363 16267 19369
rect 15979 19332 16160 19360
rect 15979 19329 15991 19332
rect 15933 19323 15991 19329
rect 15378 19252 15384 19304
rect 15436 19292 15442 19304
rect 16022 19292 16028 19304
rect 15436 19264 16028 19292
rect 15436 19252 15442 19264
rect 16022 19252 16028 19264
rect 16080 19252 16086 19304
rect 16132 19292 16160 19332
rect 16209 19329 16221 19363
rect 16255 19329 16267 19363
rect 16408 19360 16436 19459
rect 16574 19456 16580 19468
rect 16632 19456 16638 19508
rect 16758 19388 16764 19440
rect 16816 19388 16822 19440
rect 17313 19363 17371 19369
rect 17313 19360 17325 19363
rect 16209 19323 16267 19329
rect 16316 19332 16436 19360
rect 16500 19332 17325 19360
rect 16316 19292 16344 19332
rect 16132 19264 16344 19292
rect 16390 19252 16396 19304
rect 16448 19292 16454 19304
rect 16500 19292 16528 19332
rect 17313 19329 17325 19332
rect 17359 19329 17371 19363
rect 17313 19323 17371 19329
rect 16448 19264 16528 19292
rect 16448 19252 16454 19264
rect 17586 19252 17592 19304
rect 17644 19292 17650 19304
rect 25590 19292 25596 19304
rect 17644 19264 25596 19292
rect 17644 19252 17650 19264
rect 25590 19252 25596 19264
rect 25648 19252 25654 19304
rect 10928 19196 12020 19224
rect 15933 19227 15991 19233
rect 10928 19184 10934 19196
rect 15933 19193 15945 19227
rect 15979 19224 15991 19227
rect 16758 19224 16764 19236
rect 15979 19196 16764 19224
rect 15979 19193 15991 19196
rect 15933 19187 15991 19193
rect 16758 19184 16764 19196
rect 16816 19224 16822 19236
rect 16853 19227 16911 19233
rect 16853 19224 16865 19227
rect 16816 19196 16865 19224
rect 16816 19184 16822 19196
rect 16853 19193 16865 19196
rect 16899 19193 16911 19227
rect 16853 19187 16911 19193
rect 12526 19156 12532 19168
rect 7392 19128 12532 19156
rect 12526 19116 12532 19128
rect 12584 19116 12590 19168
rect 12621 19159 12679 19165
rect 12621 19125 12633 19159
rect 12667 19156 12679 19159
rect 24946 19156 24952 19168
rect 12667 19128 24952 19156
rect 12667 19125 12679 19128
rect 12621 19119 12679 19125
rect 24946 19116 24952 19128
rect 25004 19116 25010 19168
rect 1104 19066 25852 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 12214 19066
rect 12266 19014 12278 19066
rect 12330 19014 12342 19066
rect 12394 19014 12406 19066
rect 12458 19014 12470 19066
rect 12522 19014 20214 19066
rect 20266 19014 20278 19066
rect 20330 19014 20342 19066
rect 20394 19014 20406 19066
rect 20458 19014 20470 19066
rect 20522 19014 25852 19066
rect 1104 18992 25852 19014
rect 4798 18912 4804 18964
rect 4856 18912 4862 18964
rect 4890 18912 4896 18964
rect 4948 18952 4954 18964
rect 5445 18955 5503 18961
rect 5445 18952 5457 18955
rect 4948 18924 5457 18952
rect 4948 18912 4954 18924
rect 5445 18921 5457 18924
rect 5491 18921 5503 18955
rect 5445 18915 5503 18921
rect 5721 18955 5779 18961
rect 5721 18921 5733 18955
rect 5767 18952 5779 18955
rect 5810 18952 5816 18964
rect 5767 18924 5816 18952
rect 5767 18921 5779 18924
rect 5721 18915 5779 18921
rect 5810 18912 5816 18924
rect 5868 18912 5874 18964
rect 7098 18912 7104 18964
rect 7156 18912 7162 18964
rect 8570 18912 8576 18964
rect 8628 18912 8634 18964
rect 9030 18912 9036 18964
rect 9088 18912 9094 18964
rect 9401 18955 9459 18961
rect 9401 18921 9413 18955
rect 9447 18952 9459 18955
rect 9674 18952 9680 18964
rect 9447 18924 9680 18952
rect 9447 18921 9459 18924
rect 9401 18915 9459 18921
rect 9674 18912 9680 18924
rect 9732 18952 9738 18964
rect 10413 18955 10471 18961
rect 10413 18952 10425 18955
rect 9732 18924 10425 18952
rect 9732 18912 9738 18924
rect 10413 18921 10425 18924
rect 10459 18952 10471 18955
rect 10502 18952 10508 18964
rect 10459 18924 10508 18952
rect 10459 18921 10471 18924
rect 10413 18915 10471 18921
rect 10502 18912 10508 18924
rect 10560 18912 10566 18964
rect 10597 18955 10655 18961
rect 10597 18921 10609 18955
rect 10643 18952 10655 18955
rect 10870 18952 10876 18964
rect 10643 18924 10876 18952
rect 10643 18921 10655 18924
rect 10597 18915 10655 18921
rect 10870 18912 10876 18924
rect 10928 18912 10934 18964
rect 11146 18912 11152 18964
rect 11204 18952 11210 18964
rect 11882 18952 11888 18964
rect 11204 18924 11888 18952
rect 11204 18912 11210 18924
rect 11882 18912 11888 18924
rect 11940 18952 11946 18964
rect 12342 18952 12348 18964
rect 11940 18924 12348 18952
rect 11940 18912 11946 18924
rect 12342 18912 12348 18924
rect 12400 18912 12406 18964
rect 12618 18912 12624 18964
rect 12676 18952 12682 18964
rect 12713 18955 12771 18961
rect 12713 18952 12725 18955
rect 12676 18924 12725 18952
rect 12676 18912 12682 18924
rect 12713 18921 12725 18924
rect 12759 18921 12771 18955
rect 12713 18915 12771 18921
rect 14182 18912 14188 18964
rect 14240 18952 14246 18964
rect 14737 18955 14795 18961
rect 14737 18952 14749 18955
rect 14240 18924 14749 18952
rect 14240 18912 14246 18924
rect 14737 18921 14749 18924
rect 14783 18921 14795 18955
rect 14737 18915 14795 18921
rect 6822 18844 6828 18896
rect 6880 18884 6886 18896
rect 6880 18856 9536 18884
rect 6880 18844 6886 18856
rect 7742 18776 7748 18828
rect 7800 18816 7806 18828
rect 9508 18825 9536 18856
rect 10042 18844 10048 18896
rect 10100 18884 10106 18896
rect 12066 18884 12072 18896
rect 10100 18856 12072 18884
rect 10100 18844 10106 18856
rect 12066 18844 12072 18856
rect 12124 18844 12130 18896
rect 13078 18884 13084 18896
rect 12452 18856 13084 18884
rect 9493 18819 9551 18825
rect 7800 18788 8248 18816
rect 7800 18776 7806 18788
rect 3234 18708 3240 18760
rect 3292 18748 3298 18760
rect 3364 18751 3422 18757
rect 3364 18748 3376 18751
rect 3292 18720 3376 18748
rect 3292 18708 3298 18720
rect 3364 18717 3376 18720
rect 3410 18717 3422 18751
rect 3364 18711 3422 18717
rect 4433 18751 4491 18757
rect 4433 18717 4445 18751
rect 4479 18748 4491 18751
rect 4522 18748 4528 18760
rect 4479 18720 4528 18748
rect 4479 18717 4491 18720
rect 4433 18711 4491 18717
rect 4522 18708 4528 18720
rect 4580 18708 4586 18760
rect 4801 18751 4859 18757
rect 4801 18717 4813 18751
rect 4847 18748 4859 18751
rect 5261 18751 5319 18757
rect 5261 18748 5273 18751
rect 4847 18720 5273 18748
rect 4847 18717 4859 18720
rect 4801 18711 4859 18717
rect 5261 18717 5273 18720
rect 5307 18717 5319 18751
rect 5261 18711 5319 18717
rect 3467 18683 3525 18689
rect 3467 18649 3479 18683
rect 3513 18680 3525 18683
rect 3881 18683 3939 18689
rect 3881 18680 3893 18683
rect 3513 18652 3893 18680
rect 3513 18649 3525 18652
rect 3467 18643 3525 18649
rect 3881 18649 3893 18652
rect 3927 18649 3939 18683
rect 3881 18643 3939 18649
rect 3973 18683 4031 18689
rect 3973 18649 3985 18683
rect 4019 18680 4031 18683
rect 4062 18680 4068 18692
rect 4019 18652 4068 18680
rect 4019 18649 4031 18652
rect 3973 18643 4031 18649
rect 4062 18640 4068 18652
rect 4120 18680 4126 18692
rect 4816 18680 4844 18711
rect 5718 18708 5724 18760
rect 5776 18708 5782 18760
rect 5905 18751 5963 18757
rect 5905 18717 5917 18751
rect 5951 18748 5963 18751
rect 6546 18748 6552 18760
rect 5951 18720 6552 18748
rect 5951 18717 5963 18720
rect 5905 18711 5963 18717
rect 6546 18708 6552 18720
rect 6604 18708 6610 18760
rect 6914 18708 6920 18760
rect 6972 18748 6978 18760
rect 8220 18757 8248 18788
rect 9493 18785 9505 18819
rect 9539 18816 9551 18819
rect 9582 18816 9588 18828
rect 9539 18788 9588 18816
rect 9539 18785 9551 18788
rect 9493 18779 9551 18785
rect 9582 18776 9588 18788
rect 9640 18776 9646 18828
rect 10965 18819 11023 18825
rect 10965 18785 10977 18819
rect 11011 18816 11023 18819
rect 11011 18788 11442 18816
rect 11011 18785 11023 18788
rect 10965 18779 11023 18785
rect 8113 18751 8171 18757
rect 8113 18748 8125 18751
rect 6972 18720 8125 18748
rect 6972 18708 6978 18720
rect 8113 18717 8125 18720
rect 8159 18717 8171 18751
rect 8113 18711 8171 18717
rect 8205 18751 8263 18757
rect 8205 18717 8217 18751
rect 8251 18717 8263 18751
rect 8205 18711 8263 18717
rect 8389 18751 8447 18757
rect 8389 18717 8401 18751
rect 8435 18748 8447 18751
rect 9217 18751 9275 18757
rect 9217 18748 9229 18751
rect 8435 18720 9229 18748
rect 8435 18717 8447 18720
rect 8389 18711 8447 18717
rect 9217 18717 9229 18720
rect 9263 18748 9275 18751
rect 10134 18748 10140 18760
rect 9263 18720 10140 18748
rect 9263 18717 9275 18720
rect 9217 18711 9275 18717
rect 10134 18708 10140 18720
rect 10192 18708 10198 18760
rect 11238 18708 11244 18760
rect 11296 18708 11302 18760
rect 11414 18692 11442 18788
rect 11606 18776 11612 18828
rect 11664 18816 11670 18828
rect 12452 18816 12480 18856
rect 13078 18844 13084 18856
rect 13136 18844 13142 18896
rect 17586 18816 17592 18828
rect 11664 18788 12480 18816
rect 12544 18788 17592 18816
rect 11664 18776 11670 18788
rect 11514 18708 11520 18760
rect 11572 18708 11578 18760
rect 11698 18708 11704 18760
rect 11756 18708 11762 18760
rect 12161 18751 12219 18757
rect 12161 18717 12173 18751
rect 12207 18748 12219 18751
rect 12250 18748 12256 18760
rect 12207 18720 12256 18748
rect 12207 18717 12219 18720
rect 12161 18711 12219 18717
rect 12250 18708 12256 18720
rect 12308 18708 12314 18760
rect 12342 18708 12348 18760
rect 12400 18708 12406 18760
rect 12434 18708 12440 18760
rect 12492 18708 12498 18760
rect 12544 18757 12572 18788
rect 17586 18776 17592 18788
rect 17644 18776 17650 18828
rect 12529 18751 12587 18757
rect 12529 18717 12541 18751
rect 12575 18717 12587 18751
rect 12529 18711 12587 18717
rect 12618 18708 12624 18760
rect 12676 18748 12682 18760
rect 12989 18751 13047 18757
rect 12989 18748 13001 18751
rect 12676 18720 13001 18748
rect 12676 18708 12682 18720
rect 12989 18717 13001 18720
rect 13035 18717 13047 18751
rect 12989 18711 13047 18717
rect 13173 18751 13231 18757
rect 13173 18717 13185 18751
rect 13219 18748 13231 18751
rect 13354 18748 13360 18760
rect 13219 18720 13360 18748
rect 13219 18717 13231 18720
rect 13173 18711 13231 18717
rect 13354 18708 13360 18720
rect 13412 18708 13418 18760
rect 13998 18708 14004 18760
rect 14056 18748 14062 18760
rect 14185 18751 14243 18757
rect 14185 18748 14197 18751
rect 14056 18720 14197 18748
rect 14056 18708 14062 18720
rect 14185 18717 14197 18720
rect 14231 18717 14243 18751
rect 14185 18711 14243 18717
rect 14550 18708 14556 18760
rect 14608 18708 14614 18760
rect 16758 18708 16764 18760
rect 16816 18708 16822 18760
rect 17405 18751 17463 18757
rect 17405 18748 17417 18751
rect 16960 18720 17417 18748
rect 4120 18652 4844 18680
rect 7469 18683 7527 18689
rect 4120 18640 4126 18652
rect 7469 18649 7481 18683
rect 7515 18680 7527 18683
rect 7834 18680 7840 18692
rect 7515 18652 7840 18680
rect 7515 18649 7527 18652
rect 7469 18643 7527 18649
rect 7834 18640 7840 18652
rect 7892 18640 7898 18692
rect 10413 18683 10471 18689
rect 10413 18649 10425 18683
rect 10459 18680 10471 18683
rect 11146 18680 11152 18692
rect 10459 18652 11152 18680
rect 10459 18649 10471 18652
rect 10413 18643 10471 18649
rect 11146 18640 11152 18652
rect 11204 18640 11210 18692
rect 11414 18689 11428 18692
rect 11399 18683 11428 18689
rect 11399 18649 11411 18683
rect 11399 18643 11428 18649
rect 11422 18640 11428 18643
rect 11480 18640 11486 18692
rect 11609 18683 11667 18689
rect 11609 18649 11621 18683
rect 11655 18649 11667 18683
rect 11609 18643 11667 18649
rect 11885 18683 11943 18689
rect 11885 18649 11897 18683
rect 11931 18680 11943 18683
rect 13081 18683 13139 18689
rect 11931 18652 12756 18680
rect 11931 18649 11943 18652
rect 11885 18643 11943 18649
rect 4430 18572 4436 18624
rect 4488 18612 4494 18624
rect 5810 18612 5816 18624
rect 4488 18584 5816 18612
rect 4488 18572 4494 18584
rect 5810 18572 5816 18584
rect 5868 18572 5874 18624
rect 6454 18572 6460 18624
rect 6512 18612 6518 18624
rect 6733 18615 6791 18621
rect 6733 18612 6745 18615
rect 6512 18584 6745 18612
rect 6512 18572 6518 18584
rect 6733 18581 6745 18584
rect 6779 18612 6791 18615
rect 7561 18615 7619 18621
rect 7561 18612 7573 18615
rect 6779 18584 7573 18612
rect 6779 18581 6791 18584
rect 6733 18575 6791 18581
rect 7561 18581 7573 18584
rect 7607 18581 7619 18615
rect 7561 18575 7619 18581
rect 10597 18615 10655 18621
rect 10597 18581 10609 18615
rect 10643 18612 10655 18615
rect 11624 18612 11652 18643
rect 10643 18584 11652 18612
rect 12728 18612 12756 18652
rect 13081 18649 13093 18683
rect 13127 18680 13139 18683
rect 13262 18680 13268 18692
rect 13127 18652 13268 18680
rect 13127 18649 13139 18652
rect 13081 18643 13139 18649
rect 13262 18640 13268 18652
rect 13320 18680 13326 18692
rect 14369 18683 14427 18689
rect 14369 18680 14381 18683
rect 13320 18652 14381 18680
rect 13320 18640 13326 18652
rect 14369 18649 14381 18652
rect 14415 18649 14427 18683
rect 14369 18643 14427 18649
rect 14461 18683 14519 18689
rect 14461 18649 14473 18683
rect 14507 18680 14519 18683
rect 15013 18683 15071 18689
rect 15013 18680 15025 18683
rect 14507 18652 15025 18680
rect 14507 18649 14519 18652
rect 14461 18643 14519 18649
rect 15013 18649 15025 18652
rect 15059 18649 15071 18683
rect 15013 18643 15071 18649
rect 13630 18612 13636 18624
rect 12728 18584 13636 18612
rect 10643 18581 10655 18584
rect 10597 18575 10655 18581
rect 13630 18572 13636 18584
rect 13688 18572 13694 18624
rect 13814 18572 13820 18624
rect 13872 18612 13878 18624
rect 14476 18612 14504 18643
rect 15194 18640 15200 18692
rect 15252 18640 15258 18692
rect 16960 18624 16988 18720
rect 17405 18717 17417 18720
rect 17451 18717 17463 18751
rect 17405 18711 17463 18717
rect 17494 18708 17500 18760
rect 17552 18748 17558 18760
rect 17716 18751 17774 18757
rect 17716 18748 17728 18751
rect 17552 18720 17728 18748
rect 17552 18708 17558 18720
rect 17716 18717 17728 18720
rect 17762 18717 17774 18751
rect 17716 18711 17774 18717
rect 13872 18584 14504 18612
rect 13872 18572 13878 18584
rect 16942 18572 16948 18624
rect 17000 18572 17006 18624
rect 17218 18572 17224 18624
rect 17276 18572 17282 18624
rect 17819 18615 17877 18621
rect 17819 18581 17831 18615
rect 17865 18612 17877 18615
rect 18138 18612 18144 18624
rect 17865 18584 18144 18612
rect 17865 18581 17877 18584
rect 17819 18575 17877 18581
rect 18138 18572 18144 18584
rect 18196 18572 18202 18624
rect 1104 18522 25852 18544
rect 1104 18470 8214 18522
rect 8266 18470 8278 18522
rect 8330 18470 8342 18522
rect 8394 18470 8406 18522
rect 8458 18470 8470 18522
rect 8522 18470 16214 18522
rect 16266 18470 16278 18522
rect 16330 18470 16342 18522
rect 16394 18470 16406 18522
rect 16458 18470 16470 18522
rect 16522 18470 24214 18522
rect 24266 18470 24278 18522
rect 24330 18470 24342 18522
rect 24394 18470 24406 18522
rect 24458 18470 24470 18522
rect 24522 18470 25852 18522
rect 1104 18448 25852 18470
rect 3234 18368 3240 18420
rect 3292 18368 3298 18420
rect 4062 18408 4068 18420
rect 3988 18380 4068 18408
rect 3988 18349 4016 18380
rect 4062 18368 4068 18380
rect 4120 18368 4126 18420
rect 4614 18408 4620 18420
rect 4356 18380 4620 18408
rect 3973 18343 4031 18349
rect 3252 18312 3924 18340
rect 3252 18281 3280 18312
rect 3237 18275 3295 18281
rect 3237 18241 3249 18275
rect 3283 18241 3295 18275
rect 3237 18235 3295 18241
rect 3513 18275 3571 18281
rect 3513 18241 3525 18275
rect 3559 18241 3571 18275
rect 3896 18272 3924 18312
rect 3973 18309 3985 18343
rect 4019 18309 4031 18343
rect 3973 18303 4031 18309
rect 4065 18275 4123 18281
rect 4065 18272 4077 18275
rect 3896 18244 4077 18272
rect 3513 18235 3571 18241
rect 4065 18241 4077 18244
rect 4111 18272 4123 18275
rect 4246 18272 4252 18284
rect 4111 18244 4252 18272
rect 4111 18241 4123 18244
rect 4065 18235 4123 18241
rect 2869 18207 2927 18213
rect 2869 18173 2881 18207
rect 2915 18173 2927 18207
rect 3528 18204 3556 18235
rect 4246 18232 4252 18244
rect 4304 18232 4310 18284
rect 4356 18281 4384 18380
rect 4614 18368 4620 18380
rect 4672 18368 4678 18420
rect 4706 18368 4712 18420
rect 4764 18408 4770 18420
rect 5445 18411 5503 18417
rect 5445 18408 5457 18411
rect 4764 18380 5457 18408
rect 4764 18368 4770 18380
rect 5445 18377 5457 18380
rect 5491 18377 5503 18411
rect 5445 18371 5503 18377
rect 5718 18368 5724 18420
rect 5776 18408 5782 18420
rect 6457 18411 6515 18417
rect 6457 18408 6469 18411
rect 5776 18380 6469 18408
rect 5776 18368 5782 18380
rect 6457 18377 6469 18380
rect 6503 18377 6515 18411
rect 6457 18371 6515 18377
rect 6546 18368 6552 18420
rect 6604 18408 6610 18420
rect 10870 18408 10876 18420
rect 6604 18380 10876 18408
rect 6604 18368 6610 18380
rect 10870 18368 10876 18380
rect 10928 18408 10934 18420
rect 11031 18411 11089 18417
rect 11031 18408 11043 18411
rect 10928 18380 11043 18408
rect 10928 18368 10934 18380
rect 11031 18377 11043 18380
rect 11077 18377 11089 18411
rect 11031 18371 11089 18377
rect 11164 18380 11836 18408
rect 4430 18300 4436 18352
rect 4488 18300 4494 18352
rect 4632 18312 10272 18340
rect 4632 18281 4660 18312
rect 4341 18275 4399 18281
rect 4341 18241 4353 18275
rect 4387 18241 4399 18275
rect 4341 18235 4399 18241
rect 4617 18275 4675 18281
rect 4617 18241 4629 18275
rect 4663 18241 4675 18275
rect 4617 18235 4675 18241
rect 5905 18275 5963 18281
rect 5905 18241 5917 18275
rect 5951 18241 5963 18275
rect 5905 18235 5963 18241
rect 4522 18204 4528 18216
rect 3528 18176 4528 18204
rect 2869 18167 2927 18173
rect 2884 18068 2912 18167
rect 4522 18164 4528 18176
rect 4580 18204 4586 18216
rect 4801 18207 4859 18213
rect 4801 18204 4813 18207
rect 4580 18176 4813 18204
rect 4580 18164 4586 18176
rect 4801 18173 4813 18176
rect 4847 18173 4859 18207
rect 4801 18167 4859 18173
rect 5074 18164 5080 18216
rect 5132 18164 5138 18216
rect 5920 18204 5948 18235
rect 6822 18232 6828 18284
rect 6880 18232 6886 18284
rect 7469 18275 7527 18281
rect 7469 18272 7481 18275
rect 6932 18244 7481 18272
rect 5368 18176 5948 18204
rect 3237 18139 3295 18145
rect 3237 18105 3249 18139
rect 3283 18136 3295 18139
rect 4706 18136 4712 18148
rect 3283 18108 4712 18136
rect 3283 18105 3295 18108
rect 3237 18099 3295 18105
rect 4706 18096 4712 18108
rect 4764 18096 4770 18148
rect 5368 18080 5396 18176
rect 6730 18164 6736 18216
rect 6788 18204 6794 18216
rect 6932 18213 6960 18244
rect 7469 18241 7481 18244
rect 7515 18241 7527 18275
rect 7469 18235 7527 18241
rect 8941 18275 8999 18281
rect 8941 18241 8953 18275
rect 8987 18272 8999 18275
rect 9401 18275 9459 18281
rect 9401 18272 9413 18275
rect 8987 18244 9413 18272
rect 8987 18241 8999 18244
rect 8941 18235 8999 18241
rect 9401 18241 9413 18244
rect 9447 18241 9459 18275
rect 9401 18235 9459 18241
rect 9585 18275 9643 18281
rect 9585 18241 9597 18275
rect 9631 18272 9643 18275
rect 9674 18272 9680 18284
rect 9631 18244 9680 18272
rect 9631 18241 9643 18244
rect 9585 18235 9643 18241
rect 9674 18232 9680 18244
rect 9732 18232 9738 18284
rect 10244 18281 10272 18312
rect 10502 18300 10508 18352
rect 10560 18340 10566 18352
rect 11164 18340 11192 18380
rect 10560 18312 11192 18340
rect 11241 18343 11299 18349
rect 10560 18300 10566 18312
rect 11241 18309 11253 18343
rect 11287 18340 11299 18343
rect 11422 18340 11428 18352
rect 11287 18312 11428 18340
rect 11287 18309 11299 18312
rect 11241 18303 11299 18309
rect 11422 18300 11428 18312
rect 11480 18300 11486 18352
rect 11808 18340 11836 18380
rect 12250 18368 12256 18420
rect 12308 18368 12314 18420
rect 12342 18368 12348 18420
rect 12400 18408 12406 18420
rect 12529 18411 12587 18417
rect 12529 18408 12541 18411
rect 12400 18380 12541 18408
rect 12400 18368 12406 18380
rect 12529 18377 12541 18380
rect 12575 18377 12587 18411
rect 12529 18371 12587 18377
rect 12986 18368 12992 18420
rect 13044 18408 13050 18420
rect 13081 18411 13139 18417
rect 13081 18408 13093 18411
rect 13044 18380 13093 18408
rect 13044 18368 13050 18380
rect 13081 18377 13093 18380
rect 13127 18377 13139 18411
rect 13081 18371 13139 18377
rect 14185 18411 14243 18417
rect 14185 18377 14197 18411
rect 14231 18408 14243 18411
rect 15194 18408 15200 18420
rect 14231 18380 15200 18408
rect 14231 18377 14243 18380
rect 14185 18371 14243 18377
rect 13357 18343 13415 18349
rect 11808 18312 11915 18340
rect 10229 18275 10287 18281
rect 10229 18241 10241 18275
rect 10275 18241 10287 18275
rect 10229 18235 10287 18241
rect 10413 18275 10471 18281
rect 10413 18241 10425 18275
rect 10459 18272 10471 18275
rect 11514 18272 11520 18284
rect 10459 18244 11520 18272
rect 10459 18241 10471 18244
rect 10413 18235 10471 18241
rect 6917 18207 6975 18213
rect 6917 18204 6929 18207
rect 6788 18176 6929 18204
rect 6788 18164 6794 18176
rect 6917 18173 6929 18176
rect 6963 18173 6975 18207
rect 6917 18167 6975 18173
rect 7009 18207 7067 18213
rect 7009 18173 7021 18207
rect 7055 18173 7067 18207
rect 7009 18167 7067 18173
rect 9769 18207 9827 18213
rect 9769 18173 9781 18207
rect 9815 18204 9827 18207
rect 10134 18204 10140 18216
rect 9815 18176 10140 18204
rect 9815 18173 9827 18176
rect 9769 18167 9827 18173
rect 5445 18139 5503 18145
rect 5445 18105 5457 18139
rect 5491 18136 5503 18139
rect 5721 18139 5779 18145
rect 5721 18136 5733 18139
rect 5491 18108 5733 18136
rect 5491 18105 5503 18108
rect 5445 18099 5503 18105
rect 5721 18105 5733 18108
rect 5767 18105 5779 18139
rect 5721 18099 5779 18105
rect 5810 18096 5816 18148
rect 5868 18136 5874 18148
rect 7024 18136 7052 18167
rect 10134 18164 10140 18176
rect 10192 18164 10198 18216
rect 5868 18108 7052 18136
rect 9125 18139 9183 18145
rect 5868 18096 5874 18108
rect 9125 18105 9137 18139
rect 9171 18136 9183 18139
rect 9858 18136 9864 18148
rect 9171 18108 9864 18136
rect 9171 18105 9183 18108
rect 9125 18099 9183 18105
rect 9858 18096 9864 18108
rect 9916 18096 9922 18148
rect 10244 18136 10272 18235
rect 11514 18232 11520 18244
rect 11572 18232 11578 18284
rect 11606 18232 11612 18284
rect 11664 18232 11670 18284
rect 11887 18281 11915 18312
rect 13357 18309 13369 18343
rect 13403 18340 13415 18343
rect 14200 18340 14228 18371
rect 15194 18368 15200 18380
rect 15252 18408 15258 18420
rect 15289 18411 15347 18417
rect 15289 18408 15301 18411
rect 15252 18380 15301 18408
rect 15252 18368 15258 18380
rect 15289 18377 15301 18380
rect 15335 18377 15347 18411
rect 15289 18371 15347 18377
rect 15470 18368 15476 18420
rect 15528 18408 15534 18420
rect 24854 18408 24860 18420
rect 15528 18380 24860 18408
rect 15528 18368 15534 18380
rect 24854 18368 24860 18380
rect 24912 18368 24918 18420
rect 13403 18312 14228 18340
rect 13403 18309 13415 18312
rect 13357 18303 13415 18309
rect 14274 18300 14280 18352
rect 14332 18340 14338 18352
rect 16393 18343 16451 18349
rect 14332 18312 14494 18340
rect 14332 18300 14338 18312
rect 14466 18306 14494 18312
rect 16393 18309 16405 18343
rect 16439 18340 16451 18343
rect 16942 18340 16948 18352
rect 16439 18312 16948 18340
rect 16439 18309 16451 18312
rect 12066 18281 12072 18284
rect 11793 18275 11851 18281
rect 11793 18241 11805 18275
rect 11839 18241 11851 18275
rect 11793 18235 11851 18241
rect 11885 18275 11943 18281
rect 11885 18241 11897 18275
rect 11931 18241 11943 18275
rect 11885 18235 11943 18241
rect 12023 18275 12072 18281
rect 12023 18241 12035 18275
rect 12069 18241 12072 18275
rect 12023 18235 12072 18241
rect 11532 18204 11560 18232
rect 11808 18204 11836 18235
rect 12066 18232 12072 18235
rect 12124 18232 12130 18284
rect 12529 18275 12587 18281
rect 12529 18241 12541 18275
rect 12575 18241 12587 18275
rect 12529 18235 12587 18241
rect 12621 18275 12679 18281
rect 12621 18241 12633 18275
rect 12667 18272 12679 18275
rect 12710 18272 12716 18284
rect 12667 18244 12716 18272
rect 12667 18241 12679 18244
rect 12621 18235 12679 18241
rect 11532 18176 11836 18204
rect 10873 18139 10931 18145
rect 10873 18136 10885 18139
rect 10244 18108 10885 18136
rect 10873 18105 10885 18108
rect 10919 18136 10931 18139
rect 11146 18136 11152 18148
rect 10919 18108 11152 18136
rect 10919 18105 10931 18108
rect 10873 18099 10931 18105
rect 11146 18096 11152 18108
rect 11204 18096 11210 18148
rect 11330 18096 11336 18148
rect 11388 18136 11394 18148
rect 12544 18136 12572 18235
rect 12710 18232 12716 18244
rect 12768 18232 12774 18284
rect 12802 18232 12808 18284
rect 12860 18232 12866 18284
rect 13170 18232 13176 18284
rect 13228 18281 13234 18284
rect 13228 18275 13277 18281
rect 13228 18241 13231 18275
rect 13265 18241 13277 18275
rect 13228 18235 13277 18241
rect 13449 18275 13507 18281
rect 13449 18241 13461 18275
rect 13495 18241 13507 18275
rect 13630 18272 13636 18284
rect 13591 18244 13636 18272
rect 13449 18235 13507 18241
rect 13228 18232 13234 18235
rect 12618 18136 12624 18148
rect 11388 18108 12624 18136
rect 11388 18096 11394 18108
rect 12618 18096 12624 18108
rect 12676 18136 12682 18148
rect 13464 18136 13492 18235
rect 13630 18232 13636 18244
rect 13688 18232 13694 18284
rect 13722 18232 13728 18284
rect 13780 18232 13786 18284
rect 13814 18232 13820 18284
rect 13872 18272 13878 18284
rect 14466 18281 14504 18306
rect 16393 18303 16451 18309
rect 16942 18300 16948 18312
rect 17000 18340 17006 18352
rect 17000 18312 17356 18340
rect 17000 18300 17006 18312
rect 14001 18275 14059 18281
rect 14001 18272 14013 18275
rect 13872 18244 14013 18272
rect 13872 18232 13878 18244
rect 14001 18241 14013 18244
rect 14047 18241 14059 18275
rect 14001 18235 14059 18241
rect 14461 18275 14519 18281
rect 14461 18241 14473 18275
rect 14507 18241 14519 18275
rect 14461 18235 14519 18241
rect 12676 18108 13492 18136
rect 14016 18136 14044 18235
rect 14550 18232 14556 18284
rect 14608 18232 14614 18284
rect 14737 18275 14795 18281
rect 14737 18241 14749 18275
rect 14783 18241 14795 18275
rect 14737 18235 14795 18241
rect 14366 18164 14372 18216
rect 14424 18204 14430 18216
rect 14752 18204 14780 18235
rect 15194 18232 15200 18284
rect 15252 18232 15258 18284
rect 15470 18232 15476 18284
rect 15528 18232 15534 18284
rect 17328 18281 17356 18312
rect 18138 18300 18144 18352
rect 18196 18300 18202 18352
rect 15657 18275 15715 18281
rect 15657 18241 15669 18275
rect 15703 18272 15715 18275
rect 16761 18275 16819 18281
rect 16761 18272 16773 18275
rect 15703 18244 16773 18272
rect 15703 18241 15715 18244
rect 15657 18235 15715 18241
rect 16761 18241 16773 18244
rect 16807 18241 16819 18275
rect 16761 18235 16819 18241
rect 17313 18275 17371 18281
rect 17313 18241 17325 18275
rect 17359 18241 17371 18275
rect 17313 18235 17371 18241
rect 14424 18176 14780 18204
rect 14921 18207 14979 18213
rect 14424 18164 14430 18176
rect 14921 18173 14933 18207
rect 14967 18204 14979 18207
rect 15378 18204 15384 18216
rect 14967 18176 15384 18204
rect 14967 18173 14979 18176
rect 14921 18167 14979 18173
rect 15378 18164 15384 18176
rect 15436 18164 15442 18216
rect 16022 18164 16028 18216
rect 16080 18164 16086 18216
rect 16776 18204 16804 18235
rect 17589 18207 17647 18213
rect 17589 18204 17601 18207
rect 16776 18176 17601 18204
rect 17589 18173 17601 18176
rect 17635 18173 17647 18207
rect 17589 18167 17647 18173
rect 14550 18136 14556 18148
rect 14016 18108 14556 18136
rect 12676 18096 12682 18108
rect 14550 18096 14556 18108
rect 14608 18096 14614 18148
rect 17313 18139 17371 18145
rect 17313 18105 17325 18139
rect 17359 18136 17371 18139
rect 17954 18136 17960 18148
rect 17359 18108 17960 18136
rect 17359 18105 17371 18108
rect 17313 18099 17371 18105
rect 17954 18096 17960 18108
rect 18012 18136 18018 18148
rect 18049 18139 18107 18145
rect 18049 18136 18061 18139
rect 18012 18108 18061 18136
rect 18012 18096 18018 18108
rect 18049 18105 18061 18108
rect 18095 18105 18107 18139
rect 18049 18099 18107 18105
rect 4062 18068 4068 18080
rect 2884 18040 4068 18068
rect 4062 18028 4068 18040
rect 4120 18028 4126 18080
rect 4246 18028 4252 18080
rect 4304 18068 4310 18080
rect 5350 18068 5356 18080
rect 4304 18040 5356 18068
rect 4304 18028 4310 18040
rect 5350 18028 5356 18040
rect 5408 18028 5414 18080
rect 10597 18071 10655 18077
rect 10597 18037 10609 18071
rect 10643 18068 10655 18071
rect 10686 18068 10692 18080
rect 10643 18040 10692 18068
rect 10643 18037 10655 18040
rect 10597 18031 10655 18037
rect 10686 18028 10692 18040
rect 10744 18028 10750 18080
rect 11057 18071 11115 18077
rect 11057 18037 11069 18071
rect 11103 18068 11115 18071
rect 12066 18068 12072 18080
rect 11103 18040 12072 18068
rect 11103 18037 11115 18040
rect 11057 18031 11115 18037
rect 12066 18028 12072 18040
rect 12124 18028 12130 18080
rect 12710 18028 12716 18080
rect 12768 18028 12774 18080
rect 12986 18028 12992 18080
rect 13044 18068 13050 18080
rect 13354 18068 13360 18080
rect 13044 18040 13360 18068
rect 13044 18028 13050 18040
rect 13354 18028 13360 18040
rect 13412 18028 13418 18080
rect 16393 18071 16451 18077
rect 16393 18037 16405 18071
rect 16439 18068 16451 18071
rect 17494 18068 17500 18080
rect 16439 18040 17500 18068
rect 16439 18037 16451 18040
rect 16393 18031 16451 18037
rect 17494 18028 17500 18040
rect 17552 18028 17558 18080
rect 1104 17978 25852 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 12214 17978
rect 12266 17926 12278 17978
rect 12330 17926 12342 17978
rect 12394 17926 12406 17978
rect 12458 17926 12470 17978
rect 12522 17926 20214 17978
rect 20266 17926 20278 17978
rect 20330 17926 20342 17978
rect 20394 17926 20406 17978
rect 20458 17926 20470 17978
rect 20522 17926 25852 17978
rect 1104 17904 25852 17926
rect 4982 17864 4988 17876
rect 4080 17836 4988 17864
rect 4080 17737 4108 17836
rect 4982 17824 4988 17836
rect 5040 17824 5046 17876
rect 5350 17824 5356 17876
rect 5408 17824 5414 17876
rect 9033 17867 9091 17873
rect 9033 17864 9045 17867
rect 5460 17836 9045 17864
rect 4249 17799 4307 17805
rect 4249 17765 4261 17799
rect 4295 17765 4307 17799
rect 4249 17759 4307 17765
rect 4065 17731 4123 17737
rect 4065 17697 4077 17731
rect 4111 17697 4123 17731
rect 4264 17728 4292 17759
rect 4338 17756 4344 17808
rect 4396 17796 4402 17808
rect 5074 17796 5080 17808
rect 4396 17768 5080 17796
rect 4396 17756 4402 17768
rect 5074 17756 5080 17768
rect 5132 17796 5138 17808
rect 5460 17796 5488 17836
rect 9033 17833 9045 17836
rect 9079 17833 9091 17867
rect 9033 17827 9091 17833
rect 9953 17867 10011 17873
rect 9953 17833 9965 17867
rect 9999 17864 10011 17867
rect 10318 17864 10324 17876
rect 9999 17836 10324 17864
rect 9999 17833 10011 17836
rect 9953 17827 10011 17833
rect 10318 17824 10324 17836
rect 10376 17824 10382 17876
rect 11422 17864 11428 17876
rect 10520 17836 11428 17864
rect 5132 17768 5488 17796
rect 7561 17799 7619 17805
rect 5132 17756 5138 17768
rect 7561 17765 7573 17799
rect 7607 17796 7619 17799
rect 8481 17799 8539 17805
rect 8481 17796 8493 17799
rect 7607 17768 8493 17796
rect 7607 17765 7619 17768
rect 7561 17759 7619 17765
rect 8481 17765 8493 17768
rect 8527 17765 8539 17799
rect 9398 17796 9404 17808
rect 8481 17759 8539 17765
rect 9232 17768 9404 17796
rect 4264 17700 4568 17728
rect 4065 17691 4123 17697
rect 4430 17620 4436 17672
rect 4488 17620 4494 17672
rect 4540 17660 4568 17700
rect 7282 17688 7288 17740
rect 7340 17728 7346 17740
rect 7837 17731 7895 17737
rect 7837 17728 7849 17731
rect 7340 17700 7849 17728
rect 7340 17688 7346 17700
rect 7837 17697 7849 17700
rect 7883 17728 7895 17731
rect 7883 17700 8708 17728
rect 7883 17697 7895 17700
rect 7837 17691 7895 17697
rect 4706 17660 4712 17672
rect 4540 17632 4712 17660
rect 4706 17620 4712 17632
rect 4764 17660 4770 17672
rect 4826 17663 4884 17669
rect 4826 17660 4838 17663
rect 4764 17632 4838 17660
rect 4764 17620 4770 17632
rect 4826 17629 4838 17632
rect 4872 17629 4884 17663
rect 4826 17623 4884 17629
rect 5169 17663 5227 17669
rect 5169 17629 5181 17663
rect 5215 17629 5227 17663
rect 5169 17623 5227 17629
rect 4338 17552 4344 17604
rect 4396 17592 4402 17604
rect 5184 17592 5212 17623
rect 5626 17620 5632 17672
rect 5684 17620 5690 17672
rect 5721 17663 5779 17669
rect 5721 17629 5733 17663
rect 5767 17660 5779 17663
rect 5810 17660 5816 17672
rect 5767 17632 5816 17660
rect 5767 17629 5779 17632
rect 5721 17623 5779 17629
rect 5810 17620 5816 17632
rect 5868 17620 5874 17672
rect 5905 17663 5963 17669
rect 5905 17629 5917 17663
rect 5951 17660 5963 17663
rect 6546 17660 6552 17672
rect 5951 17632 6552 17660
rect 5951 17629 5963 17632
rect 5905 17623 5963 17629
rect 6546 17620 6552 17632
rect 6604 17620 6610 17672
rect 6917 17663 6975 17669
rect 6917 17629 6929 17663
rect 6963 17660 6975 17663
rect 7006 17660 7012 17672
rect 6963 17632 7012 17660
rect 6963 17629 6975 17632
rect 6917 17623 6975 17629
rect 7006 17620 7012 17632
rect 7064 17620 7070 17672
rect 7193 17663 7251 17669
rect 7193 17629 7205 17663
rect 7239 17660 7251 17663
rect 8205 17663 8263 17669
rect 8205 17660 8217 17663
rect 7239 17632 8217 17660
rect 7239 17629 7251 17632
rect 7193 17623 7251 17629
rect 8205 17629 8217 17632
rect 8251 17660 8263 17663
rect 8570 17660 8576 17672
rect 8251 17632 8576 17660
rect 8251 17629 8263 17632
rect 8205 17623 8263 17629
rect 8570 17620 8576 17632
rect 8628 17620 8634 17672
rect 8680 17669 8708 17700
rect 9232 17669 9260 17768
rect 9398 17756 9404 17768
rect 9456 17796 9462 17808
rect 9769 17799 9827 17805
rect 9769 17796 9781 17799
rect 9456 17768 9781 17796
rect 9456 17756 9462 17768
rect 9769 17765 9781 17768
rect 9815 17765 9827 17799
rect 10520 17796 10548 17836
rect 11422 17824 11428 17836
rect 11480 17824 11486 17876
rect 11514 17824 11520 17876
rect 11572 17824 11578 17876
rect 11882 17824 11888 17876
rect 11940 17864 11946 17876
rect 11977 17867 12035 17873
rect 11977 17864 11989 17867
rect 11940 17836 11989 17864
rect 11940 17824 11946 17836
rect 11977 17833 11989 17836
rect 12023 17833 12035 17867
rect 12986 17864 12992 17876
rect 11977 17827 12035 17833
rect 12406 17836 12992 17864
rect 9769 17759 9827 17765
rect 10336 17768 10548 17796
rect 10226 17728 10232 17740
rect 9416 17700 10232 17728
rect 9416 17669 9444 17700
rect 10226 17688 10232 17700
rect 10284 17688 10290 17740
rect 8665 17663 8723 17669
rect 8665 17629 8677 17663
rect 8711 17629 8723 17663
rect 8665 17623 8723 17629
rect 9217 17663 9275 17669
rect 9217 17629 9229 17663
rect 9263 17629 9275 17663
rect 9217 17623 9275 17629
rect 9401 17663 9459 17669
rect 9401 17629 9413 17663
rect 9447 17629 9459 17663
rect 9401 17623 9459 17629
rect 9493 17663 9551 17669
rect 9493 17629 9505 17663
rect 9539 17660 9551 17663
rect 9766 17660 9772 17672
rect 9539 17632 9772 17660
rect 9539 17629 9551 17632
rect 9493 17623 9551 17629
rect 9766 17620 9772 17632
rect 9824 17620 9830 17672
rect 10336 17660 10364 17768
rect 10594 17756 10600 17808
rect 10652 17796 10658 17808
rect 12406 17796 12434 17836
rect 12986 17824 12992 17836
rect 13044 17824 13050 17876
rect 13078 17824 13084 17876
rect 13136 17864 13142 17876
rect 13725 17867 13783 17873
rect 13725 17864 13737 17867
rect 13136 17836 13737 17864
rect 13136 17824 13142 17836
rect 13725 17833 13737 17836
rect 13771 17833 13783 17867
rect 13725 17827 13783 17833
rect 15381 17867 15439 17873
rect 15381 17833 15393 17867
rect 15427 17864 15439 17867
rect 15562 17864 15568 17876
rect 15427 17836 15568 17864
rect 15427 17833 15439 17836
rect 15381 17827 15439 17833
rect 10652 17768 12434 17796
rect 12529 17799 12587 17805
rect 10652 17756 10658 17768
rect 12529 17765 12541 17799
rect 12575 17796 12587 17799
rect 12710 17796 12716 17808
rect 12575 17768 12716 17796
rect 12575 17765 12587 17768
rect 12529 17759 12587 17765
rect 12710 17756 12716 17768
rect 12768 17756 12774 17808
rect 12802 17756 12808 17808
rect 12860 17796 12866 17808
rect 13262 17796 13268 17808
rect 12860 17768 13268 17796
rect 12860 17756 12866 17768
rect 13262 17756 13268 17768
rect 13320 17756 13326 17808
rect 13740 17796 13768 17827
rect 15562 17824 15568 17836
rect 15620 17824 15626 17876
rect 15933 17867 15991 17873
rect 15933 17833 15945 17867
rect 15979 17864 15991 17867
rect 16022 17864 16028 17876
rect 15979 17836 16028 17864
rect 15979 17833 15991 17836
rect 15933 17827 15991 17833
rect 16022 17824 16028 17836
rect 16080 17824 16086 17876
rect 15470 17796 15476 17808
rect 13740 17768 15476 17796
rect 15470 17756 15476 17768
rect 15528 17756 15534 17808
rect 17037 17799 17095 17805
rect 17037 17765 17049 17799
rect 17083 17796 17095 17799
rect 17218 17796 17224 17808
rect 17083 17768 17224 17796
rect 17083 17765 17095 17768
rect 17037 17759 17095 17765
rect 17218 17756 17224 17768
rect 17276 17756 17282 17808
rect 10505 17731 10563 17737
rect 10505 17697 10517 17731
rect 10551 17728 10563 17731
rect 13814 17728 13820 17740
rect 10551 17700 12388 17728
rect 10551 17697 10563 17700
rect 10505 17691 10563 17697
rect 9952 17635 10364 17660
rect 9907 17632 10364 17635
rect 9907 17629 9980 17632
rect 4396 17564 5212 17592
rect 9907 17595 9919 17629
rect 9953 17598 9980 17629
rect 10410 17620 10416 17672
rect 10468 17620 10474 17672
rect 10594 17620 10600 17672
rect 10652 17620 10658 17672
rect 10873 17663 10931 17669
rect 10873 17629 10885 17663
rect 10919 17660 10931 17663
rect 10962 17660 10968 17672
rect 10919 17632 10968 17660
rect 10919 17629 10931 17632
rect 10873 17623 10931 17629
rect 10962 17620 10968 17632
rect 11020 17620 11026 17672
rect 11057 17663 11115 17669
rect 11057 17629 11069 17663
rect 11103 17629 11115 17663
rect 12161 17663 12219 17669
rect 12161 17660 12173 17663
rect 11057 17623 11115 17629
rect 11564 17632 12173 17660
rect 9953 17595 9965 17598
rect 9907 17589 9965 17595
rect 4396 17552 4402 17564
rect 10134 17552 10140 17604
rect 10192 17552 10198 17604
rect 10778 17592 10784 17604
rect 10428 17564 10784 17592
rect 4430 17484 4436 17536
rect 4488 17524 4494 17536
rect 4755 17527 4813 17533
rect 4755 17524 4767 17527
rect 4488 17496 4767 17524
rect 4488 17484 4494 17496
rect 4755 17493 4767 17496
rect 4801 17493 4813 17527
rect 4755 17487 4813 17493
rect 5810 17484 5816 17536
rect 5868 17524 5874 17536
rect 6089 17527 6147 17533
rect 6089 17524 6101 17527
rect 5868 17496 6101 17524
rect 5868 17484 5874 17496
rect 6089 17493 6101 17496
rect 6135 17493 6147 17527
rect 6089 17487 6147 17493
rect 6178 17484 6184 17536
rect 6236 17524 6242 17536
rect 6733 17527 6791 17533
rect 6733 17524 6745 17527
rect 6236 17496 6745 17524
rect 6236 17484 6242 17496
rect 6733 17493 6745 17496
rect 6779 17493 6791 17527
rect 6733 17487 6791 17493
rect 7558 17484 7564 17536
rect 7616 17524 7622 17536
rect 7837 17527 7895 17533
rect 7837 17524 7849 17527
rect 7616 17496 7849 17524
rect 7616 17484 7622 17496
rect 7837 17493 7849 17496
rect 7883 17493 7895 17527
rect 7837 17487 7895 17493
rect 7926 17484 7932 17536
rect 7984 17524 7990 17536
rect 10428 17524 10456 17564
rect 10778 17552 10784 17564
rect 10836 17592 10842 17604
rect 11072 17592 11100 17623
rect 10836 17564 11100 17592
rect 10836 17552 10842 17564
rect 11146 17552 11152 17604
rect 11204 17592 11210 17604
rect 11564 17601 11592 17632
rect 12161 17629 12173 17632
rect 12207 17629 12219 17663
rect 12161 17623 12219 17629
rect 12253 17663 12311 17669
rect 12253 17629 12265 17663
rect 12299 17660 12311 17663
rect 12360 17660 12388 17700
rect 12820 17700 13820 17728
rect 12299 17632 12388 17660
rect 12299 17629 12311 17632
rect 12253 17623 12311 17629
rect 12710 17620 12716 17672
rect 12768 17660 12774 17672
rect 12820 17669 12848 17700
rect 13814 17688 13820 17700
rect 13872 17688 13878 17740
rect 15933 17731 15991 17737
rect 15933 17697 15945 17731
rect 15979 17728 15991 17731
rect 16669 17731 16727 17737
rect 16669 17728 16681 17731
rect 15979 17700 16681 17728
rect 15979 17697 15991 17700
rect 15933 17691 15991 17697
rect 16669 17697 16681 17700
rect 16715 17697 16727 17731
rect 16669 17691 16727 17697
rect 12805 17663 12863 17669
rect 12805 17660 12817 17663
rect 12768 17632 12817 17660
rect 12768 17620 12774 17632
rect 12805 17629 12817 17632
rect 12851 17629 12863 17663
rect 12805 17623 12863 17629
rect 12986 17620 12992 17672
rect 13044 17620 13050 17672
rect 13446 17620 13452 17672
rect 13504 17620 13510 17672
rect 13630 17620 13636 17672
rect 13688 17660 13694 17672
rect 14185 17663 14243 17669
rect 14185 17660 14197 17663
rect 13688 17632 14197 17660
rect 13688 17620 13694 17632
rect 14185 17629 14197 17632
rect 14231 17629 14243 17663
rect 14185 17623 14243 17629
rect 14278 17663 14336 17669
rect 14278 17629 14290 17663
rect 14324 17660 14336 17663
rect 14366 17660 14372 17672
rect 14324 17632 14372 17660
rect 14324 17629 14336 17632
rect 14278 17623 14336 17629
rect 11333 17595 11391 17601
rect 11333 17592 11345 17595
rect 11204 17564 11345 17592
rect 11204 17552 11210 17564
rect 11333 17561 11345 17564
rect 11379 17561 11391 17595
rect 11333 17555 11391 17561
rect 11549 17595 11607 17601
rect 11549 17561 11561 17595
rect 11595 17561 11607 17595
rect 11549 17555 11607 17561
rect 13725 17595 13783 17601
rect 13725 17561 13737 17595
rect 13771 17561 13783 17595
rect 13725 17555 13783 17561
rect 7984 17496 10456 17524
rect 7984 17484 7990 17496
rect 10870 17484 10876 17536
rect 10928 17484 10934 17536
rect 11701 17527 11759 17533
rect 11701 17493 11713 17527
rect 11747 17524 11759 17527
rect 11790 17524 11796 17536
rect 11747 17496 11796 17524
rect 11747 17493 11759 17496
rect 11701 17487 11759 17493
rect 11790 17484 11796 17496
rect 11848 17484 11854 17536
rect 12158 17484 12164 17536
rect 12216 17484 12222 17536
rect 12250 17484 12256 17536
rect 12308 17524 12314 17536
rect 12345 17527 12403 17533
rect 12345 17524 12357 17527
rect 12308 17496 12357 17524
rect 12308 17484 12314 17496
rect 12345 17493 12357 17496
rect 12391 17524 12403 17527
rect 12802 17524 12808 17536
rect 12391 17496 12808 17524
rect 12391 17493 12403 17496
rect 12345 17487 12403 17493
rect 12802 17484 12808 17496
rect 12860 17484 12866 17536
rect 12894 17484 12900 17536
rect 12952 17484 12958 17536
rect 12986 17484 12992 17536
rect 13044 17524 13050 17536
rect 13541 17527 13599 17533
rect 13541 17524 13553 17527
rect 13044 17496 13553 17524
rect 13044 17484 13050 17496
rect 13541 17493 13553 17496
rect 13587 17493 13599 17527
rect 13740 17524 13768 17555
rect 13814 17552 13820 17604
rect 13872 17592 13878 17604
rect 14292 17592 14320 17623
rect 14366 17620 14372 17632
rect 14424 17620 14430 17672
rect 14642 17620 14648 17672
rect 14700 17669 14706 17672
rect 14700 17660 14708 17669
rect 14700 17632 14745 17660
rect 14700 17623 14708 17632
rect 14700 17620 14706 17623
rect 15562 17620 15568 17672
rect 15620 17620 15626 17672
rect 16022 17620 16028 17672
rect 16080 17660 16086 17672
rect 16117 17663 16175 17669
rect 16117 17660 16129 17663
rect 16080 17632 16129 17660
rect 16080 17620 16086 17632
rect 16117 17629 16129 17632
rect 16163 17629 16175 17663
rect 16117 17623 16175 17629
rect 16393 17663 16451 17669
rect 16393 17629 16405 17663
rect 16439 17629 16451 17663
rect 16393 17623 16451 17629
rect 13872 17564 14320 17592
rect 13872 17552 13878 17564
rect 14458 17552 14464 17604
rect 14516 17552 14522 17604
rect 14553 17595 14611 17601
rect 14553 17561 14565 17595
rect 14599 17561 14611 17595
rect 14553 17555 14611 17561
rect 13906 17524 13912 17536
rect 13740 17496 13912 17524
rect 13541 17487 13599 17493
rect 13906 17484 13912 17496
rect 13964 17524 13970 17536
rect 14274 17524 14280 17536
rect 13964 17496 14280 17524
rect 13964 17484 13970 17496
rect 14274 17484 14280 17496
rect 14332 17524 14338 17536
rect 14568 17524 14596 17555
rect 15930 17552 15936 17604
rect 15988 17592 15994 17604
rect 16408 17592 16436 17623
rect 17954 17620 17960 17672
rect 18012 17620 18018 17672
rect 18601 17663 18659 17669
rect 18601 17660 18613 17663
rect 18248 17632 18613 17660
rect 18248 17604 18276 17632
rect 18601 17629 18613 17632
rect 18647 17629 18659 17663
rect 18601 17623 18659 17629
rect 15988 17564 16436 17592
rect 18141 17595 18199 17601
rect 15988 17552 15994 17564
rect 18141 17561 18153 17595
rect 18187 17592 18199 17595
rect 18230 17592 18236 17604
rect 18187 17564 18236 17592
rect 18187 17561 18199 17564
rect 18141 17555 18199 17561
rect 18230 17552 18236 17564
rect 18288 17552 18294 17604
rect 14332 17496 14596 17524
rect 14332 17484 14338 17496
rect 14826 17484 14832 17536
rect 14884 17484 14890 17536
rect 16114 17484 16120 17536
rect 16172 17524 16178 17536
rect 16301 17527 16359 17533
rect 16301 17524 16313 17527
rect 16172 17496 16313 17524
rect 16172 17484 16178 17496
rect 16301 17493 16313 17496
rect 16347 17493 16359 17527
rect 16301 17487 16359 17493
rect 17037 17527 17095 17533
rect 17037 17493 17049 17527
rect 17083 17524 17095 17527
rect 17494 17524 17500 17536
rect 17083 17496 17500 17524
rect 17083 17493 17095 17496
rect 17037 17487 17095 17493
rect 17494 17484 17500 17496
rect 17552 17484 17558 17536
rect 18414 17484 18420 17536
rect 18472 17484 18478 17536
rect 1104 17434 25852 17456
rect 1104 17382 8214 17434
rect 8266 17382 8278 17434
rect 8330 17382 8342 17434
rect 8394 17382 8406 17434
rect 8458 17382 8470 17434
rect 8522 17382 16214 17434
rect 16266 17382 16278 17434
rect 16330 17382 16342 17434
rect 16394 17382 16406 17434
rect 16458 17382 16470 17434
rect 16522 17382 24214 17434
rect 24266 17382 24278 17434
rect 24330 17382 24342 17434
rect 24394 17382 24406 17434
rect 24458 17382 24470 17434
rect 24522 17382 25852 17434
rect 1104 17360 25852 17382
rect 4706 17280 4712 17332
rect 4764 17280 4770 17332
rect 8849 17323 8907 17329
rect 8849 17320 8861 17323
rect 5368 17292 8861 17320
rect 3513 17255 3571 17261
rect 3513 17221 3525 17255
rect 3559 17252 3571 17255
rect 4338 17252 4344 17264
rect 3559 17224 4344 17252
rect 3559 17221 3571 17224
rect 3513 17215 3571 17221
rect 4338 17212 4344 17224
rect 4396 17212 4402 17264
rect 4430 17212 4436 17264
rect 4488 17212 4494 17264
rect 4522 17212 4528 17264
rect 4580 17252 4586 17264
rect 5368 17252 5396 17292
rect 8849 17289 8861 17292
rect 8895 17289 8907 17323
rect 10870 17320 10876 17332
rect 8849 17283 8907 17289
rect 9232 17292 10876 17320
rect 4580 17224 5396 17252
rect 4580 17212 4586 17224
rect 3053 17187 3111 17193
rect 3053 17153 3065 17187
rect 3099 17153 3111 17187
rect 3053 17147 3111 17153
rect 3605 17187 3663 17193
rect 3605 17153 3617 17187
rect 3651 17184 3663 17187
rect 4982 17184 4988 17196
rect 3651 17156 4988 17184
rect 3651 17153 3663 17156
rect 3605 17147 3663 17153
rect 3068 17116 3096 17147
rect 4982 17144 4988 17156
rect 5040 17144 5046 17196
rect 5092 17193 5120 17224
rect 7006 17212 7012 17264
rect 7064 17212 7070 17264
rect 5077 17187 5135 17193
rect 5077 17153 5089 17187
rect 5123 17153 5135 17187
rect 5077 17147 5135 17153
rect 5353 17187 5411 17193
rect 5353 17153 5365 17187
rect 5399 17184 5411 17187
rect 5810 17184 5816 17196
rect 5399 17156 5816 17184
rect 5399 17153 5411 17156
rect 5353 17147 5411 17153
rect 5810 17144 5816 17156
rect 5868 17144 5874 17196
rect 5905 17187 5963 17193
rect 5905 17153 5917 17187
rect 5951 17184 5963 17187
rect 6086 17184 6092 17196
rect 5951 17156 6092 17184
rect 5951 17153 5963 17156
rect 5905 17147 5963 17153
rect 6086 17144 6092 17156
rect 6144 17144 6150 17196
rect 6508 17187 6566 17193
rect 6508 17153 6520 17187
rect 6554 17184 6566 17187
rect 7558 17184 7564 17196
rect 6554 17156 7564 17184
rect 6554 17153 6566 17156
rect 6508 17147 6566 17153
rect 7558 17144 7564 17156
rect 7616 17144 7622 17196
rect 7926 17144 7932 17196
rect 7984 17144 7990 17196
rect 8113 17187 8171 17193
rect 8113 17153 8125 17187
rect 8159 17184 8171 17187
rect 8386 17184 8392 17196
rect 8159 17156 8392 17184
rect 8159 17153 8171 17156
rect 8113 17147 8171 17153
rect 8386 17144 8392 17156
rect 8444 17144 8450 17196
rect 8573 17187 8631 17193
rect 8573 17153 8585 17187
rect 8619 17153 8631 17187
rect 8573 17147 8631 17153
rect 9033 17187 9091 17193
rect 9033 17153 9045 17187
rect 9079 17153 9091 17187
rect 9033 17147 9091 17153
rect 3878 17116 3884 17128
rect 3068 17088 3884 17116
rect 3878 17076 3884 17088
rect 3936 17076 3942 17128
rect 4706 17076 4712 17128
rect 4764 17076 4770 17128
rect 6595 17119 6653 17125
rect 6595 17085 6607 17119
rect 6641 17116 6653 17119
rect 6917 17119 6975 17125
rect 6917 17116 6929 17119
rect 6641 17088 6929 17116
rect 6641 17085 6653 17088
rect 6595 17079 6653 17085
rect 6917 17085 6929 17088
rect 6963 17085 6975 17119
rect 6917 17079 6975 17085
rect 7466 17076 7472 17128
rect 7524 17076 7530 17128
rect 8021 17119 8079 17125
rect 8021 17085 8033 17119
rect 8067 17116 8079 17119
rect 8478 17116 8484 17128
rect 8067 17088 8484 17116
rect 8067 17085 8079 17088
rect 8021 17079 8079 17085
rect 8478 17076 8484 17088
rect 8536 17076 8542 17128
rect 5902 16940 5908 16992
rect 5960 16940 5966 16992
rect 7834 16940 7840 16992
rect 7892 16980 7898 16992
rect 8481 16983 8539 16989
rect 8481 16980 8493 16983
rect 7892 16952 8493 16980
rect 7892 16940 7898 16952
rect 8481 16949 8493 16952
rect 8527 16949 8539 16983
rect 8588 16980 8616 17147
rect 9048 17116 9076 17147
rect 9122 17144 9128 17196
rect 9180 17144 9186 17196
rect 9232 17193 9260 17292
rect 10870 17280 10876 17292
rect 10928 17320 10934 17332
rect 11977 17323 12035 17329
rect 11977 17320 11989 17323
rect 10928 17292 11989 17320
rect 10928 17280 10934 17292
rect 11977 17289 11989 17292
rect 12023 17289 12035 17323
rect 11977 17283 12035 17289
rect 12158 17280 12164 17332
rect 12216 17320 12222 17332
rect 12529 17323 12587 17329
rect 12529 17320 12541 17323
rect 12216 17292 12541 17320
rect 12216 17280 12222 17292
rect 12529 17289 12541 17292
rect 12575 17289 12587 17323
rect 12529 17283 12587 17289
rect 12894 17280 12900 17332
rect 12952 17320 12958 17332
rect 13998 17320 14004 17332
rect 12952 17292 14004 17320
rect 12952 17280 12958 17292
rect 13998 17280 14004 17292
rect 14056 17280 14062 17332
rect 14090 17280 14096 17332
rect 14148 17320 14154 17332
rect 14148 17292 14412 17320
rect 14148 17280 14154 17292
rect 10060 17224 13032 17252
rect 9217 17187 9275 17193
rect 9217 17153 9229 17187
rect 9263 17153 9275 17187
rect 9217 17147 9275 17153
rect 9398 17144 9404 17196
rect 9456 17144 9462 17196
rect 9674 17144 9680 17196
rect 9732 17144 9738 17196
rect 9858 17144 9864 17196
rect 9916 17144 9922 17196
rect 9950 17144 9956 17196
rect 10008 17144 10014 17196
rect 10060 17193 10088 17224
rect 10045 17187 10103 17193
rect 10045 17153 10057 17187
rect 10091 17153 10103 17187
rect 10045 17147 10103 17153
rect 10134 17144 10140 17196
rect 10192 17184 10198 17196
rect 10502 17184 10508 17196
rect 10192 17156 10508 17184
rect 10192 17144 10198 17156
rect 10502 17144 10508 17156
rect 10560 17144 10566 17196
rect 10594 17144 10600 17196
rect 10652 17144 10658 17196
rect 11057 17187 11115 17193
rect 11057 17153 11069 17187
rect 11103 17184 11115 17187
rect 11238 17184 11244 17196
rect 11103 17156 11244 17184
rect 11103 17153 11115 17156
rect 11057 17147 11115 17153
rect 11238 17144 11244 17156
rect 11296 17144 11302 17196
rect 11422 17144 11428 17196
rect 11480 17184 11486 17196
rect 11885 17187 11943 17193
rect 11480 17183 11560 17184
rect 11624 17183 11744 17184
rect 11885 17183 11897 17187
rect 11480 17156 11897 17183
rect 11480 17144 11486 17156
rect 11532 17155 11652 17156
rect 11716 17155 11897 17156
rect 11885 17153 11897 17155
rect 11931 17153 11943 17187
rect 11885 17147 11943 17153
rect 12618 17144 12624 17196
rect 12676 17184 12682 17196
rect 12713 17187 12771 17193
rect 12713 17184 12725 17187
rect 12676 17156 12725 17184
rect 12676 17144 12682 17156
rect 12713 17153 12725 17156
rect 12759 17153 12771 17187
rect 12713 17147 12771 17153
rect 12802 17144 12808 17196
rect 12860 17144 12866 17196
rect 12894 17144 12900 17196
rect 12952 17144 12958 17196
rect 13004 17184 13032 17224
rect 13004 17156 13400 17184
rect 11768 17119 11826 17125
rect 9048 17088 11008 17116
rect 10980 17060 11008 17088
rect 11768 17085 11780 17119
rect 11814 17116 11826 17119
rect 11814 17108 11915 17116
rect 11814 17088 11928 17108
rect 11814 17085 11826 17088
rect 11768 17079 11826 17085
rect 11887 17080 11928 17088
rect 9122 17008 9128 17060
rect 9180 17048 9186 17060
rect 9490 17048 9496 17060
rect 9180 17020 9496 17048
rect 9180 17008 9186 17020
rect 9490 17008 9496 17020
rect 9548 17048 9554 17060
rect 9950 17048 9956 17060
rect 9548 17020 9956 17048
rect 9548 17008 9554 17020
rect 9950 17008 9956 17020
rect 10008 17048 10014 17060
rect 10008 17020 10180 17048
rect 10008 17008 10014 17020
rect 10042 16980 10048 16992
rect 8588 16952 10048 16980
rect 8481 16943 8539 16949
rect 10042 16940 10048 16952
rect 10100 16940 10106 16992
rect 10152 16980 10180 17020
rect 10226 17008 10232 17060
rect 10284 17008 10290 17060
rect 10962 17008 10968 17060
rect 11020 17008 11026 17060
rect 11149 17051 11207 17057
rect 11149 17017 11161 17051
rect 11195 17048 11207 17051
rect 11330 17048 11336 17060
rect 11195 17020 11336 17048
rect 11195 17017 11207 17020
rect 11149 17011 11207 17017
rect 11330 17008 11336 17020
rect 11388 17008 11394 17060
rect 11606 17008 11612 17060
rect 11664 17008 11670 17060
rect 11900 17048 11928 17080
rect 12066 17076 12072 17128
rect 12124 17116 12130 17128
rect 12253 17119 12311 17125
rect 12253 17116 12265 17119
rect 12124 17088 12265 17116
rect 12124 17076 12130 17088
rect 12253 17085 12265 17088
rect 12299 17085 12311 17119
rect 12253 17079 12311 17085
rect 13262 17076 13268 17128
rect 13320 17076 13326 17128
rect 13372 17116 13400 17156
rect 13446 17144 13452 17196
rect 13504 17144 13510 17196
rect 13541 17187 13599 17193
rect 13541 17153 13553 17187
rect 13587 17184 13599 17187
rect 13722 17184 13728 17196
rect 13587 17156 13728 17184
rect 13587 17153 13599 17156
rect 13541 17147 13599 17153
rect 13722 17144 13728 17156
rect 13780 17144 13786 17196
rect 14016 17193 14044 17280
rect 14274 17212 14280 17264
rect 14332 17212 14338 17264
rect 14001 17187 14059 17193
rect 14001 17153 14013 17187
rect 14047 17153 14059 17187
rect 14001 17147 14059 17153
rect 14182 17144 14188 17196
rect 14240 17144 14246 17196
rect 14384 17193 14412 17292
rect 14826 17212 14832 17264
rect 14884 17252 14890 17264
rect 14884 17224 20760 17252
rect 14884 17212 14890 17224
rect 16942 17193 16948 17196
rect 14369 17187 14427 17193
rect 14369 17153 14381 17187
rect 14415 17153 14427 17187
rect 14369 17147 14427 17153
rect 16910 17187 16948 17193
rect 16910 17153 16922 17187
rect 16910 17147 16948 17153
rect 16942 17144 16948 17147
rect 17000 17144 17006 17196
rect 17328 17193 17356 17224
rect 17313 17187 17371 17193
rect 17313 17153 17325 17187
rect 17359 17153 17371 17187
rect 17313 17147 17371 17153
rect 18230 17144 18236 17196
rect 18288 17144 18294 17196
rect 19334 17144 19340 17196
rect 19392 17144 19398 17196
rect 20732 17193 20760 17224
rect 20717 17187 20775 17193
rect 20717 17153 20729 17187
rect 20763 17153 20775 17187
rect 20717 17147 20775 17153
rect 18877 17119 18935 17125
rect 13372 17088 18736 17116
rect 11974 17048 11980 17060
rect 11900 17020 11980 17048
rect 11974 17008 11980 17020
rect 12032 17008 12038 17060
rect 12158 17008 12164 17060
rect 12216 17048 12222 17060
rect 13357 17051 13415 17057
rect 13357 17048 13369 17051
rect 12216 17020 13369 17048
rect 12216 17008 12222 17020
rect 13357 17017 13369 17020
rect 13403 17017 13415 17051
rect 13357 17011 13415 17017
rect 17126 17008 17132 17060
rect 17184 17048 17190 17060
rect 18601 17051 18659 17057
rect 18601 17048 18613 17051
rect 17184 17020 18613 17048
rect 17184 17008 17190 17020
rect 18601 17017 18613 17020
rect 18647 17017 18659 17051
rect 18708 17048 18736 17088
rect 18877 17085 18889 17119
rect 18923 17116 18935 17119
rect 19245 17119 19303 17125
rect 19245 17116 19257 17119
rect 18923 17088 19257 17116
rect 18923 17085 18935 17088
rect 18877 17079 18935 17085
rect 19245 17085 19257 17088
rect 19291 17085 19303 17119
rect 19245 17079 19303 17085
rect 19518 17048 19524 17060
rect 18708 17020 19524 17048
rect 18601 17011 18659 17017
rect 19518 17008 19524 17020
rect 19576 17008 19582 17060
rect 10689 16983 10747 16989
rect 10689 16980 10701 16983
rect 10152 16952 10701 16980
rect 10689 16949 10701 16952
rect 10735 16949 10747 16983
rect 10689 16943 10747 16949
rect 14550 16940 14556 16992
rect 14608 16940 14614 16992
rect 16574 16940 16580 16992
rect 16632 16980 16638 16992
rect 16807 16983 16865 16989
rect 16807 16980 16819 16983
rect 16632 16952 16819 16980
rect 16632 16940 16638 16952
rect 16807 16949 16819 16952
rect 16853 16949 16865 16983
rect 16807 16943 16865 16949
rect 17034 16940 17040 16992
rect 17092 16980 17098 16992
rect 21542 16980 21548 16992
rect 17092 16952 21548 16980
rect 17092 16940 17098 16952
rect 21542 16940 21548 16952
rect 21600 16940 21606 16992
rect 1104 16890 25852 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 12214 16890
rect 12266 16838 12278 16890
rect 12330 16838 12342 16890
rect 12394 16838 12406 16890
rect 12458 16838 12470 16890
rect 12522 16838 20214 16890
rect 20266 16838 20278 16890
rect 20330 16838 20342 16890
rect 20394 16838 20406 16890
rect 20458 16838 20470 16890
rect 20522 16838 25852 16890
rect 1104 16816 25852 16838
rect 3878 16736 3884 16788
rect 3936 16776 3942 16788
rect 4433 16779 4491 16785
rect 4433 16776 4445 16779
rect 3936 16748 4445 16776
rect 3936 16736 3942 16748
rect 4433 16745 4445 16748
rect 4479 16745 4491 16779
rect 4433 16739 4491 16745
rect 4706 16736 4712 16788
rect 4764 16776 4770 16788
rect 4801 16779 4859 16785
rect 4801 16776 4813 16779
rect 4764 16748 4813 16776
rect 4764 16736 4770 16748
rect 4801 16745 4813 16748
rect 4847 16745 4859 16779
rect 4801 16739 4859 16745
rect 7006 16736 7012 16788
rect 7064 16776 7070 16788
rect 7101 16779 7159 16785
rect 7101 16776 7113 16779
rect 7064 16748 7113 16776
rect 7064 16736 7070 16748
rect 7101 16745 7113 16748
rect 7147 16745 7159 16779
rect 7101 16739 7159 16745
rect 8570 16736 8576 16788
rect 8628 16776 8634 16788
rect 9585 16779 9643 16785
rect 9585 16776 9597 16779
rect 8628 16748 9597 16776
rect 8628 16736 8634 16748
rect 9585 16745 9597 16748
rect 9631 16745 9643 16779
rect 9585 16739 9643 16745
rect 11149 16779 11207 16785
rect 11149 16745 11161 16779
rect 11195 16776 11207 16779
rect 11514 16776 11520 16788
rect 11195 16748 11520 16776
rect 11195 16745 11207 16748
rect 11149 16739 11207 16745
rect 11514 16736 11520 16748
rect 11572 16736 11578 16788
rect 11606 16736 11612 16788
rect 11664 16736 11670 16788
rect 11882 16736 11888 16788
rect 11940 16776 11946 16788
rect 23566 16776 23572 16788
rect 11940 16748 23572 16776
rect 11940 16736 11946 16748
rect 23566 16736 23572 16748
rect 23624 16736 23630 16788
rect 5261 16711 5319 16717
rect 5261 16677 5273 16711
rect 5307 16677 5319 16711
rect 5261 16671 5319 16677
rect 3970 16532 3976 16584
rect 4028 16532 4034 16584
rect 4246 16532 4252 16584
rect 4304 16532 4310 16584
rect 4982 16532 4988 16584
rect 5040 16572 5046 16584
rect 5276 16572 5304 16671
rect 5902 16668 5908 16720
rect 5960 16708 5966 16720
rect 6181 16711 6239 16717
rect 6181 16708 6193 16711
rect 5960 16680 6193 16708
rect 5960 16668 5966 16680
rect 6181 16677 6193 16680
rect 6227 16677 6239 16711
rect 10597 16711 10655 16717
rect 6181 16671 6239 16677
rect 8680 16680 10548 16708
rect 5920 16640 5948 16668
rect 7466 16640 7472 16652
rect 5644 16612 5948 16640
rect 7024 16612 7472 16640
rect 5040 16544 5304 16572
rect 5445 16575 5503 16581
rect 5040 16532 5046 16544
rect 5445 16541 5457 16575
rect 5491 16572 5503 16575
rect 5644 16572 5672 16612
rect 5491 16544 5672 16572
rect 5721 16575 5779 16581
rect 5491 16541 5503 16544
rect 5445 16535 5503 16541
rect 5721 16541 5733 16575
rect 5767 16572 5779 16575
rect 5810 16572 5816 16584
rect 5767 16544 5816 16572
rect 5767 16541 5779 16544
rect 5721 16535 5779 16541
rect 5810 16532 5816 16544
rect 5868 16532 5874 16584
rect 6549 16575 6607 16581
rect 6549 16541 6561 16575
rect 6595 16572 6607 16575
rect 7024 16572 7052 16612
rect 7466 16600 7472 16612
rect 7524 16640 7530 16652
rect 7837 16643 7895 16649
rect 7837 16640 7849 16643
rect 7524 16612 7849 16640
rect 7524 16600 7530 16612
rect 7837 16609 7849 16612
rect 7883 16609 7895 16643
rect 7837 16603 7895 16609
rect 6595 16544 7052 16572
rect 7101 16575 7159 16581
rect 6595 16541 6607 16544
rect 6549 16535 6607 16541
rect 7101 16541 7113 16575
rect 7147 16572 7159 16575
rect 7282 16572 7288 16584
rect 7147 16544 7288 16572
rect 7147 16541 7159 16544
rect 7101 16535 7159 16541
rect 7282 16532 7288 16544
rect 7340 16532 7346 16584
rect 7374 16532 7380 16584
rect 7432 16532 7438 16584
rect 7650 16532 7656 16584
rect 7708 16532 7714 16584
rect 8386 16532 8392 16584
rect 8444 16572 8450 16584
rect 8680 16581 8708 16680
rect 9306 16640 9312 16652
rect 9232 16612 9312 16640
rect 8481 16575 8539 16581
rect 8481 16572 8493 16575
rect 8444 16544 8493 16572
rect 8444 16532 8450 16544
rect 8481 16541 8493 16544
rect 8527 16541 8539 16575
rect 8481 16535 8539 16541
rect 8665 16575 8723 16581
rect 8665 16541 8677 16575
rect 8711 16541 8723 16575
rect 8665 16535 8723 16541
rect 6270 16464 6276 16516
rect 6328 16464 6334 16516
rect 7469 16507 7527 16513
rect 7469 16473 7481 16507
rect 7515 16504 7527 16507
rect 7742 16504 7748 16516
rect 7515 16476 7748 16504
rect 7515 16473 7527 16476
rect 7469 16467 7527 16473
rect 7742 16464 7748 16476
rect 7800 16464 7806 16516
rect 8496 16504 8524 16535
rect 8754 16532 8760 16584
rect 8812 16572 8818 16584
rect 9232 16581 9260 16612
rect 9306 16600 9312 16612
rect 9364 16600 9370 16652
rect 9582 16600 9588 16652
rect 9640 16640 9646 16652
rect 9640 16612 9904 16640
rect 9640 16600 9646 16612
rect 9876 16581 9904 16612
rect 10520 16584 10548 16680
rect 10597 16677 10609 16711
rect 10643 16708 10655 16711
rect 11974 16708 11980 16720
rect 10643 16680 11980 16708
rect 10643 16677 10655 16680
rect 10597 16671 10655 16677
rect 11974 16668 11980 16680
rect 12032 16708 12038 16720
rect 12250 16708 12256 16720
rect 12032 16680 12256 16708
rect 12032 16668 12038 16680
rect 12250 16668 12256 16680
rect 12308 16668 12314 16720
rect 12618 16708 12624 16720
rect 12544 16680 12624 16708
rect 11606 16640 11612 16652
rect 11256 16612 11612 16640
rect 9033 16575 9091 16581
rect 9033 16572 9045 16575
rect 8812 16544 9045 16572
rect 8812 16532 8818 16544
rect 9033 16541 9045 16544
rect 9079 16541 9091 16575
rect 9033 16535 9091 16541
rect 9217 16575 9275 16581
rect 9217 16541 9229 16575
rect 9263 16541 9275 16575
rect 9217 16535 9275 16541
rect 9401 16575 9459 16581
rect 9401 16541 9413 16575
rect 9447 16572 9459 16575
rect 9861 16575 9919 16581
rect 9447 16544 9812 16572
rect 9447 16541 9459 16544
rect 9401 16535 9459 16541
rect 8846 16504 8852 16516
rect 8496 16476 8852 16504
rect 8846 16464 8852 16476
rect 8904 16464 8910 16516
rect 9122 16464 9128 16516
rect 9180 16504 9186 16516
rect 9309 16507 9367 16513
rect 9309 16504 9321 16507
rect 9180 16476 9321 16504
rect 9180 16464 9186 16476
rect 9309 16473 9321 16476
rect 9355 16473 9367 16507
rect 9674 16504 9680 16516
rect 9309 16467 9367 16473
rect 9416 16476 9680 16504
rect 4065 16439 4123 16445
rect 4065 16405 4077 16439
rect 4111 16436 4123 16439
rect 4154 16436 4160 16448
rect 4111 16408 4160 16436
rect 4111 16405 4123 16408
rect 4065 16399 4123 16405
rect 4154 16396 4160 16408
rect 4212 16436 4218 16448
rect 5718 16436 5724 16448
rect 4212 16408 5724 16436
rect 4212 16396 4218 16408
rect 5718 16396 5724 16408
rect 5776 16396 5782 16448
rect 8665 16439 8723 16445
rect 8665 16405 8677 16439
rect 8711 16436 8723 16439
rect 9416 16436 9444 16476
rect 9674 16464 9680 16476
rect 9732 16464 9738 16516
rect 9784 16504 9812 16544
rect 9861 16541 9873 16575
rect 9907 16541 9919 16575
rect 9861 16535 9919 16541
rect 10134 16532 10140 16584
rect 10192 16532 10198 16584
rect 10502 16532 10508 16584
rect 10560 16532 10566 16584
rect 10689 16575 10747 16581
rect 10689 16541 10701 16575
rect 10735 16572 10747 16575
rect 10870 16572 10876 16584
rect 10735 16544 10876 16572
rect 10735 16541 10747 16544
rect 10689 16535 10747 16541
rect 10870 16532 10876 16544
rect 10928 16532 10934 16584
rect 11256 16581 11284 16612
rect 11606 16600 11612 16612
rect 11664 16600 11670 16652
rect 12544 16640 12572 16680
rect 12618 16668 12624 16680
rect 12676 16708 12682 16720
rect 12802 16708 12808 16720
rect 12676 16680 12808 16708
rect 12676 16668 12682 16680
rect 12802 16668 12808 16680
rect 12860 16668 12866 16720
rect 12986 16668 12992 16720
rect 13044 16708 13050 16720
rect 13449 16711 13507 16717
rect 13449 16708 13461 16711
rect 13044 16680 13461 16708
rect 13044 16668 13050 16680
rect 13449 16677 13461 16680
rect 13495 16677 13507 16711
rect 13449 16671 13507 16677
rect 14461 16711 14519 16717
rect 14461 16677 14473 16711
rect 14507 16708 14519 16711
rect 14918 16708 14924 16720
rect 14507 16680 14924 16708
rect 14507 16677 14519 16680
rect 14461 16671 14519 16677
rect 14918 16668 14924 16680
rect 14976 16668 14982 16720
rect 16022 16668 16028 16720
rect 16080 16668 16086 16720
rect 16485 16711 16543 16717
rect 16485 16677 16497 16711
rect 16531 16708 16543 16711
rect 16531 16680 16896 16708
rect 16531 16677 16543 16680
rect 16485 16671 16543 16677
rect 12084 16612 12572 16640
rect 12728 16612 13124 16640
rect 11240 16575 11298 16581
rect 11240 16541 11252 16575
rect 11286 16541 11298 16575
rect 11240 16535 11298 16541
rect 11330 16532 11336 16584
rect 11388 16532 11394 16584
rect 11514 16532 11520 16584
rect 11572 16572 11578 16584
rect 11793 16575 11851 16581
rect 11793 16572 11805 16575
rect 11572 16544 11805 16572
rect 11572 16532 11578 16544
rect 11793 16541 11805 16544
rect 11839 16541 11851 16575
rect 11793 16535 11851 16541
rect 11977 16575 12035 16581
rect 11977 16541 11989 16575
rect 12023 16572 12035 16575
rect 12084 16572 12112 16612
rect 12023 16544 12112 16572
rect 12023 16541 12035 16544
rect 11977 16535 12035 16541
rect 12158 16532 12164 16584
rect 12216 16532 12222 16584
rect 12526 16532 12532 16584
rect 12584 16572 12590 16584
rect 12728 16581 12756 16612
rect 12712 16575 12770 16581
rect 12584 16566 12664 16572
rect 12712 16566 12724 16575
rect 12584 16544 12724 16566
rect 12584 16532 12590 16544
rect 12636 16541 12724 16544
rect 12758 16541 12770 16575
rect 12636 16538 12770 16541
rect 12712 16535 12770 16538
rect 12802 16532 12808 16584
rect 12860 16532 12866 16584
rect 13096 16581 13124 16612
rect 13538 16600 13544 16652
rect 13596 16640 13602 16652
rect 16040 16640 16068 16668
rect 13596 16612 13860 16640
rect 13596 16600 13602 16612
rect 13081 16575 13139 16581
rect 13081 16541 13093 16575
rect 13127 16541 13139 16575
rect 13081 16535 13139 16541
rect 13170 16532 13176 16584
rect 13228 16572 13234 16584
rect 13265 16575 13323 16581
rect 13265 16572 13277 16575
rect 13228 16544 13277 16572
rect 13228 16532 13234 16544
rect 13265 16541 13277 16544
rect 13311 16572 13323 16575
rect 13722 16572 13728 16584
rect 13311 16544 13728 16572
rect 13311 16541 13323 16544
rect 13265 16535 13323 16541
rect 13722 16532 13728 16544
rect 13780 16532 13786 16584
rect 13832 16572 13860 16612
rect 14936 16612 16160 16640
rect 14737 16575 14795 16581
rect 14737 16572 14749 16575
rect 13832 16544 14749 16572
rect 14737 16541 14749 16544
rect 14783 16572 14795 16575
rect 14936 16572 14964 16612
rect 14783 16544 14964 16572
rect 14783 16541 14795 16544
rect 14737 16535 14795 16541
rect 15102 16532 15108 16584
rect 15160 16532 15166 16584
rect 15746 16532 15752 16584
rect 15804 16572 15810 16584
rect 16132 16581 16160 16612
rect 16758 16600 16764 16652
rect 16816 16600 16822 16652
rect 16868 16640 16896 16680
rect 16942 16668 16948 16720
rect 17000 16668 17006 16720
rect 18414 16668 18420 16720
rect 18472 16668 18478 16720
rect 17405 16643 17463 16649
rect 17405 16640 17417 16643
rect 16868 16612 17417 16640
rect 17405 16609 17417 16612
rect 17451 16640 17463 16643
rect 18049 16643 18107 16649
rect 18049 16640 18061 16643
rect 17451 16612 18061 16640
rect 17451 16609 17463 16612
rect 17405 16603 17463 16609
rect 18049 16609 18061 16612
rect 18095 16609 18107 16643
rect 18049 16603 18107 16609
rect 15933 16575 15991 16581
rect 15933 16572 15945 16575
rect 15804 16544 15945 16572
rect 15804 16532 15810 16544
rect 15933 16541 15945 16544
rect 15979 16541 15991 16575
rect 15933 16535 15991 16541
rect 16117 16575 16175 16581
rect 16117 16541 16129 16575
rect 16163 16541 16175 16575
rect 16117 16535 16175 16541
rect 16206 16532 16212 16584
rect 16264 16532 16270 16584
rect 16301 16575 16359 16581
rect 16301 16541 16313 16575
rect 16347 16572 16359 16575
rect 17773 16575 17831 16581
rect 16347 16544 17724 16572
rect 16347 16541 16359 16544
rect 16301 16535 16359 16541
rect 11885 16507 11943 16513
rect 9784 16476 11836 16504
rect 11808 16448 11836 16476
rect 11885 16473 11897 16507
rect 11931 16504 11943 16507
rect 12066 16504 12072 16516
rect 11931 16476 12072 16504
rect 11931 16473 11943 16476
rect 11885 16467 11943 16473
rect 12066 16464 12072 16476
rect 12124 16464 12130 16516
rect 12250 16464 12256 16516
rect 12308 16504 12314 16516
rect 14921 16507 14979 16513
rect 14921 16504 14933 16507
rect 12308 16476 14933 16504
rect 12308 16464 12314 16476
rect 14921 16473 14933 16476
rect 14967 16473 14979 16507
rect 14921 16467 14979 16473
rect 15013 16507 15071 16513
rect 15013 16473 15025 16507
rect 15059 16504 15071 16507
rect 15378 16504 15384 16516
rect 15059 16476 15384 16504
rect 15059 16473 15071 16476
rect 15013 16467 15071 16473
rect 15378 16464 15384 16476
rect 15436 16464 15442 16516
rect 15657 16507 15715 16513
rect 15657 16473 15669 16507
rect 15703 16504 15715 16507
rect 16316 16504 16344 16535
rect 15703 16476 16344 16504
rect 15703 16473 15715 16476
rect 15657 16467 15715 16473
rect 17126 16464 17132 16516
rect 17184 16464 17190 16516
rect 17696 16504 17724 16544
rect 17773 16541 17785 16575
rect 17819 16572 17831 16575
rect 18230 16572 18236 16584
rect 17819 16544 18236 16572
rect 17819 16541 17831 16544
rect 17773 16535 17831 16541
rect 18230 16532 18236 16544
rect 18288 16532 18294 16584
rect 18877 16575 18935 16581
rect 18877 16541 18889 16575
rect 18923 16572 18935 16575
rect 19334 16572 19340 16584
rect 18923 16544 19340 16572
rect 18923 16541 18935 16544
rect 18877 16535 18935 16541
rect 19334 16532 19340 16544
rect 19392 16532 19398 16584
rect 26142 16504 26148 16516
rect 17696 16476 26148 16504
rect 26142 16464 26148 16476
rect 26200 16464 26206 16516
rect 8711 16408 9444 16436
rect 8711 16405 8723 16408
rect 8665 16399 8723 16405
rect 9490 16396 9496 16448
rect 9548 16436 9554 16448
rect 10137 16439 10195 16445
rect 10137 16436 10149 16439
rect 9548 16408 10149 16436
rect 9548 16396 9554 16408
rect 10137 16405 10149 16408
rect 10183 16436 10195 16439
rect 11238 16436 11244 16448
rect 10183 16408 11244 16436
rect 10183 16405 10195 16408
rect 10137 16399 10195 16405
rect 11238 16396 11244 16408
rect 11296 16396 11302 16448
rect 11790 16396 11796 16448
rect 11848 16396 11854 16448
rect 12434 16396 12440 16448
rect 12492 16396 12498 16448
rect 15289 16439 15347 16445
rect 15289 16405 15301 16439
rect 15335 16436 15347 16439
rect 16758 16436 16764 16448
rect 15335 16408 16764 16436
rect 15335 16405 15347 16408
rect 15289 16399 15347 16405
rect 16758 16396 16764 16408
rect 16816 16396 16822 16448
rect 17773 16439 17831 16445
rect 17773 16405 17785 16439
rect 17819 16436 17831 16439
rect 18417 16439 18475 16445
rect 18417 16436 18429 16439
rect 17819 16408 18429 16436
rect 17819 16405 17831 16408
rect 17773 16399 17831 16405
rect 18417 16405 18429 16408
rect 18463 16436 18475 16439
rect 18693 16439 18751 16445
rect 18693 16436 18705 16439
rect 18463 16408 18705 16436
rect 18463 16405 18475 16408
rect 18417 16399 18475 16405
rect 18693 16405 18705 16408
rect 18739 16405 18751 16439
rect 18693 16399 18751 16405
rect 1104 16346 25852 16368
rect 1104 16294 8214 16346
rect 8266 16294 8278 16346
rect 8330 16294 8342 16346
rect 8394 16294 8406 16346
rect 8458 16294 8470 16346
rect 8522 16294 16214 16346
rect 16266 16294 16278 16346
rect 16330 16294 16342 16346
rect 16394 16294 16406 16346
rect 16458 16294 16470 16346
rect 16522 16294 24214 16346
rect 24266 16294 24278 16346
rect 24330 16294 24342 16346
rect 24394 16294 24406 16346
rect 24458 16294 24470 16346
rect 24522 16294 25852 16346
rect 1104 16272 25852 16294
rect 6089 16235 6147 16241
rect 6089 16201 6101 16235
rect 6135 16232 6147 16235
rect 6825 16235 6883 16241
rect 6825 16232 6837 16235
rect 6135 16204 6837 16232
rect 6135 16201 6147 16204
rect 6089 16195 6147 16201
rect 6825 16201 6837 16204
rect 6871 16201 6883 16235
rect 6825 16195 6883 16201
rect 7650 16192 7656 16244
rect 7708 16232 7714 16244
rect 8757 16235 8815 16241
rect 8757 16232 8769 16235
rect 7708 16204 8769 16232
rect 7708 16192 7714 16204
rect 8757 16201 8769 16204
rect 8803 16201 8815 16235
rect 8757 16195 8815 16201
rect 8846 16192 8852 16244
rect 8904 16232 8910 16244
rect 9490 16232 9496 16244
rect 8904 16204 9496 16232
rect 8904 16192 8910 16204
rect 9490 16192 9496 16204
rect 9548 16192 9554 16244
rect 10778 16192 10784 16244
rect 10836 16232 10842 16244
rect 10873 16235 10931 16241
rect 10873 16232 10885 16235
rect 10836 16204 10885 16232
rect 10836 16192 10842 16204
rect 10873 16201 10885 16204
rect 10919 16201 10931 16235
rect 10873 16195 10931 16201
rect 11606 16192 11612 16244
rect 11664 16192 11670 16244
rect 11790 16192 11796 16244
rect 11848 16232 11854 16244
rect 12986 16232 12992 16244
rect 11848 16204 12992 16232
rect 11848 16192 11854 16204
rect 12986 16192 12992 16204
rect 13044 16192 13050 16244
rect 13081 16235 13139 16241
rect 13081 16201 13093 16235
rect 13127 16232 13139 16235
rect 13262 16232 13268 16244
rect 13127 16204 13268 16232
rect 13127 16201 13139 16204
rect 13081 16195 13139 16201
rect 13262 16192 13268 16204
rect 13320 16192 13326 16244
rect 13354 16192 13360 16244
rect 13412 16192 13418 16244
rect 14182 16192 14188 16244
rect 14240 16192 14246 16244
rect 15102 16192 15108 16244
rect 15160 16232 15166 16244
rect 15160 16204 16344 16232
rect 15160 16192 15166 16204
rect 4246 16124 4252 16176
rect 4304 16164 4310 16176
rect 9677 16167 9735 16173
rect 9677 16164 9689 16167
rect 4304 16136 9689 16164
rect 4304 16124 4310 16136
rect 9677 16133 9689 16136
rect 9723 16133 9735 16167
rect 9677 16127 9735 16133
rect 10502 16124 10508 16176
rect 10560 16164 10566 16176
rect 11974 16164 11980 16176
rect 10560 16136 11980 16164
rect 10560 16124 10566 16136
rect 11974 16124 11980 16136
rect 12032 16164 12038 16176
rect 12526 16164 12532 16176
rect 12032 16136 12532 16164
rect 12032 16124 12038 16136
rect 12526 16124 12532 16136
rect 12584 16164 12590 16176
rect 13372 16164 13400 16192
rect 12584 16136 12664 16164
rect 13372 16136 14412 16164
rect 12584 16124 12590 16136
rect 3237 16099 3295 16105
rect 3237 16065 3249 16099
rect 3283 16065 3295 16099
rect 3237 16059 3295 16065
rect 3050 15988 3056 16040
rect 3108 16028 3114 16040
rect 3252 16028 3280 16059
rect 3418 16056 3424 16108
rect 3476 16096 3482 16108
rect 4154 16096 4160 16108
rect 3476 16068 4160 16096
rect 3476 16056 3482 16068
rect 4154 16056 4160 16068
rect 4212 16056 4218 16108
rect 4341 16099 4399 16105
rect 4341 16065 4353 16099
rect 4387 16065 4399 16099
rect 4341 16059 4399 16065
rect 4356 16028 4384 16059
rect 6086 16056 6092 16108
rect 6144 16096 6150 16108
rect 7285 16099 7343 16105
rect 7285 16096 7297 16099
rect 6144 16068 7297 16096
rect 6144 16056 6150 16068
rect 7285 16065 7297 16068
rect 7331 16065 7343 16099
rect 7285 16059 7343 16065
rect 7745 16099 7803 16105
rect 7745 16065 7757 16099
rect 7791 16096 7803 16099
rect 8294 16096 8300 16108
rect 7791 16068 8300 16096
rect 7791 16065 7803 16068
rect 7745 16059 7803 16065
rect 8294 16056 8300 16068
rect 8352 16056 8358 16108
rect 8941 16099 8999 16105
rect 8941 16065 8953 16099
rect 8987 16096 8999 16099
rect 9122 16096 9128 16108
rect 8987 16068 9128 16096
rect 8987 16065 8999 16068
rect 8941 16059 8999 16065
rect 9122 16056 9128 16068
rect 9180 16056 9186 16108
rect 9214 16056 9220 16108
rect 9272 16056 9278 16108
rect 9306 16056 9312 16108
rect 9364 16096 9370 16108
rect 9401 16099 9459 16105
rect 9401 16096 9413 16099
rect 9364 16068 9413 16096
rect 9364 16056 9370 16068
rect 9401 16065 9413 16068
rect 9447 16096 9459 16099
rect 9861 16099 9919 16105
rect 9861 16096 9873 16099
rect 9447 16068 9873 16096
rect 9447 16065 9459 16068
rect 9401 16059 9459 16065
rect 9861 16065 9873 16068
rect 9907 16065 9919 16099
rect 9861 16059 9919 16065
rect 10137 16099 10195 16105
rect 10137 16065 10149 16099
rect 10183 16096 10195 16099
rect 10686 16096 10692 16108
rect 10183 16068 10692 16096
rect 10183 16065 10195 16068
rect 10137 16059 10195 16065
rect 10686 16056 10692 16068
rect 10744 16056 10750 16108
rect 11057 16099 11115 16105
rect 11057 16065 11069 16099
rect 11103 16065 11115 16099
rect 11057 16059 11115 16065
rect 11241 16099 11299 16105
rect 11241 16065 11253 16099
rect 11287 16096 11299 16099
rect 11330 16096 11336 16108
rect 11287 16068 11336 16096
rect 11287 16065 11299 16068
rect 11241 16059 11299 16065
rect 3108 16000 4384 16028
rect 3108 15988 3114 16000
rect 4356 15960 4384 16000
rect 5721 16031 5779 16037
rect 5721 15997 5733 16031
rect 5767 16028 5779 16031
rect 6457 16031 6515 16037
rect 6457 16028 6469 16031
rect 5767 16000 6469 16028
rect 5767 15997 5779 16000
rect 5721 15991 5779 15997
rect 6457 15997 6469 16000
rect 6503 16028 6515 16031
rect 10226 16028 10232 16040
rect 6503 16000 10232 16028
rect 6503 15997 6515 16000
rect 6457 15991 6515 15997
rect 10226 15988 10232 16000
rect 10284 15988 10290 16040
rect 6825 15963 6883 15969
rect 4356 15932 6224 15960
rect 3142 15852 3148 15904
rect 3200 15892 3206 15904
rect 3237 15895 3295 15901
rect 3237 15892 3249 15895
rect 3200 15864 3249 15892
rect 3200 15852 3206 15864
rect 3237 15861 3249 15864
rect 3283 15861 3295 15895
rect 3237 15855 3295 15861
rect 4341 15895 4399 15901
rect 4341 15861 4353 15895
rect 4387 15892 4399 15895
rect 4614 15892 4620 15904
rect 4387 15864 4620 15892
rect 4387 15861 4399 15864
rect 4341 15855 4399 15861
rect 4614 15852 4620 15864
rect 4672 15852 4678 15904
rect 6086 15852 6092 15904
rect 6144 15852 6150 15904
rect 6196 15892 6224 15932
rect 6825 15929 6837 15963
rect 6871 15960 6883 15963
rect 7101 15963 7159 15969
rect 7101 15960 7113 15963
rect 6871 15932 7113 15960
rect 6871 15929 6883 15932
rect 6825 15923 6883 15929
rect 7101 15929 7113 15932
rect 7147 15929 7159 15963
rect 7101 15923 7159 15929
rect 7742 15920 7748 15972
rect 7800 15960 7806 15972
rect 7929 15963 7987 15969
rect 7929 15960 7941 15963
rect 7800 15932 7941 15960
rect 7800 15920 7806 15932
rect 7929 15929 7941 15932
rect 7975 15929 7987 15963
rect 7929 15923 7987 15929
rect 9582 15920 9588 15972
rect 9640 15960 9646 15972
rect 9953 15963 10011 15969
rect 9953 15960 9965 15963
rect 9640 15932 9965 15960
rect 9640 15920 9646 15932
rect 9953 15929 9965 15932
rect 9999 15929 10011 15963
rect 9953 15923 10011 15929
rect 10042 15920 10048 15972
rect 10100 15920 10106 15972
rect 11072 15960 11100 16059
rect 11330 16056 11336 16068
rect 11388 16056 11394 16108
rect 11422 16056 11428 16108
rect 11480 16096 11486 16108
rect 11793 16099 11851 16105
rect 11793 16096 11805 16099
rect 11480 16068 11805 16096
rect 11480 16056 11486 16068
rect 11793 16065 11805 16068
rect 11839 16065 11851 16099
rect 11793 16059 11851 16065
rect 11885 16099 11943 16105
rect 11885 16065 11897 16099
rect 11931 16065 11943 16099
rect 11885 16059 11943 16065
rect 12161 16099 12219 16105
rect 12161 16065 12173 16099
rect 12207 16096 12219 16099
rect 12434 16096 12440 16108
rect 12207 16068 12440 16096
rect 12207 16065 12219 16068
rect 12161 16059 12219 16065
rect 11146 15988 11152 16040
rect 11204 16028 11210 16040
rect 11900 16028 11928 16059
rect 12434 16056 12440 16068
rect 12492 16056 12498 16108
rect 12636 16105 12664 16136
rect 12621 16099 12679 16105
rect 12621 16065 12633 16099
rect 12667 16065 12679 16099
rect 12621 16059 12679 16065
rect 12710 16056 12716 16108
rect 12768 16056 12774 16108
rect 12802 16056 12808 16108
rect 12860 16096 12866 16108
rect 14384 16105 14412 16136
rect 14550 16124 14556 16176
rect 14608 16164 14614 16176
rect 14829 16167 14887 16173
rect 14829 16164 14841 16167
rect 14608 16136 14841 16164
rect 14608 16124 14614 16136
rect 14829 16133 14841 16136
rect 14875 16133 14887 16167
rect 14829 16127 14887 16133
rect 15562 16124 15568 16176
rect 15620 16164 15626 16176
rect 16117 16167 16175 16173
rect 16117 16164 16129 16167
rect 15620 16136 16129 16164
rect 15620 16124 15626 16136
rect 16117 16133 16129 16136
rect 16163 16164 16175 16167
rect 16206 16164 16212 16176
rect 16163 16136 16212 16164
rect 16163 16133 16175 16136
rect 16117 16127 16175 16133
rect 16206 16124 16212 16136
rect 16264 16124 16270 16176
rect 14185 16099 14243 16105
rect 14185 16096 14197 16099
rect 12860 16068 14197 16096
rect 12860 16056 12866 16068
rect 14185 16065 14197 16068
rect 14231 16065 14243 16099
rect 14185 16059 14243 16065
rect 14369 16099 14427 16105
rect 14369 16065 14381 16099
rect 14415 16065 14427 16099
rect 14369 16059 14427 16065
rect 15013 16099 15071 16105
rect 15013 16065 15025 16099
rect 15059 16096 15071 16099
rect 15102 16096 15108 16108
rect 15059 16068 15108 16096
rect 15059 16065 15071 16068
rect 15013 16059 15071 16065
rect 15102 16056 15108 16068
rect 15160 16056 15166 16108
rect 15197 16099 15255 16105
rect 15197 16065 15209 16099
rect 15243 16096 15255 16099
rect 15473 16099 15531 16105
rect 15473 16096 15485 16099
rect 15243 16068 15485 16096
rect 15243 16065 15255 16068
rect 15197 16059 15255 16065
rect 15473 16065 15485 16068
rect 15519 16065 15531 16099
rect 15473 16059 15531 16065
rect 11204 16000 11928 16028
rect 11204 15988 11210 16000
rect 12066 15988 12072 16040
rect 12124 15988 12130 16040
rect 12894 16028 12900 16040
rect 12406 16000 12900 16028
rect 11514 15960 11520 15972
rect 11072 15932 11520 15960
rect 11514 15920 11520 15932
rect 11572 15960 11578 15972
rect 12406 15960 12434 16000
rect 12894 15988 12900 16000
rect 12952 16028 12958 16040
rect 12952 16000 13492 16028
rect 12952 15988 12958 16000
rect 13464 15969 13492 16000
rect 13722 15988 13728 16040
rect 13780 16028 13786 16040
rect 13817 16031 13875 16037
rect 13817 16028 13829 16031
rect 13780 16000 13829 16028
rect 13780 15988 13786 16000
rect 13817 15997 13829 16000
rect 13863 15997 13875 16031
rect 16316 16028 16344 16204
rect 16942 16192 16948 16244
rect 17000 16232 17006 16244
rect 17129 16235 17187 16241
rect 17129 16232 17141 16235
rect 17000 16204 17141 16232
rect 17000 16192 17006 16204
rect 17129 16201 17141 16204
rect 17175 16201 17187 16235
rect 17129 16195 17187 16201
rect 16393 16167 16451 16173
rect 16393 16133 16405 16167
rect 16439 16164 16451 16167
rect 16439 16136 17172 16164
rect 16439 16133 16451 16136
rect 16393 16127 16451 16133
rect 17144 16108 17172 16136
rect 16758 16056 16764 16108
rect 16816 16056 16822 16108
rect 17126 16056 17132 16108
rect 17184 16096 17190 16108
rect 17589 16099 17647 16105
rect 17589 16096 17601 16099
rect 17184 16068 17601 16096
rect 17184 16056 17190 16068
rect 17589 16065 17601 16068
rect 17635 16065 17647 16099
rect 17589 16059 17647 16065
rect 26418 16028 26424 16040
rect 16316 16000 26424 16028
rect 13817 15991 13875 15997
rect 26418 15988 26424 16000
rect 26476 15988 26482 16040
rect 11572 15932 12434 15960
rect 13449 15963 13507 15969
rect 11572 15920 11578 15932
rect 13449 15929 13461 15963
rect 13495 15929 13507 15963
rect 13449 15923 13507 15929
rect 17129 15963 17187 15969
rect 17129 15929 17141 15963
rect 17175 15960 17187 15963
rect 17405 15963 17463 15969
rect 17405 15960 17417 15963
rect 17175 15932 17417 15960
rect 17175 15929 17187 15932
rect 17129 15923 17187 15929
rect 17405 15929 17417 15932
rect 17451 15929 17463 15963
rect 17405 15923 17463 15929
rect 8018 15892 8024 15904
rect 6196 15864 8024 15892
rect 8018 15852 8024 15864
rect 8076 15892 8082 15904
rect 9858 15892 9864 15904
rect 8076 15864 9864 15892
rect 8076 15852 8082 15864
rect 9858 15852 9864 15864
rect 9916 15852 9922 15904
rect 10318 15852 10324 15904
rect 10376 15892 10382 15904
rect 11698 15892 11704 15904
rect 10376 15864 11704 15892
rect 10376 15852 10382 15864
rect 11698 15852 11704 15864
rect 11756 15852 11762 15904
rect 12986 15852 12992 15904
rect 13044 15892 13050 15904
rect 17310 15892 17316 15904
rect 13044 15864 17316 15892
rect 13044 15852 13050 15864
rect 17310 15852 17316 15864
rect 17368 15852 17374 15904
rect 1104 15802 25852 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 12214 15802
rect 12266 15750 12278 15802
rect 12330 15750 12342 15802
rect 12394 15750 12406 15802
rect 12458 15750 12470 15802
rect 12522 15750 20214 15802
rect 20266 15750 20278 15802
rect 20330 15750 20342 15802
rect 20394 15750 20406 15802
rect 20458 15750 20470 15802
rect 20522 15750 25852 15802
rect 1104 15728 25852 15750
rect 3418 15688 3424 15700
rect 2608 15660 3424 15688
rect 2501 15487 2559 15493
rect 2501 15453 2513 15487
rect 2547 15484 2559 15487
rect 2608 15484 2636 15660
rect 3418 15648 3424 15660
rect 3476 15648 3482 15700
rect 6270 15648 6276 15700
rect 6328 15688 6334 15700
rect 6411 15691 6469 15697
rect 6411 15688 6423 15691
rect 6328 15660 6423 15688
rect 6328 15648 6334 15660
rect 6411 15657 6423 15660
rect 6457 15657 6469 15691
rect 6411 15651 6469 15657
rect 8665 15691 8723 15697
rect 8665 15657 8677 15691
rect 8711 15657 8723 15691
rect 8665 15651 8723 15657
rect 3050 15620 3056 15632
rect 2700 15592 3056 15620
rect 2700 15493 2728 15592
rect 3050 15580 3056 15592
rect 3108 15580 3114 15632
rect 5718 15580 5724 15632
rect 5776 15620 5782 15632
rect 7009 15623 7067 15629
rect 7009 15620 7021 15623
rect 5776 15592 7021 15620
rect 5776 15580 5782 15592
rect 7009 15589 7021 15592
rect 7055 15589 7067 15623
rect 8680 15620 8708 15651
rect 9214 15648 9220 15700
rect 9272 15688 9278 15700
rect 9272 15660 10548 15688
rect 9272 15648 9278 15660
rect 8680 15592 9628 15620
rect 7009 15583 7067 15589
rect 3234 15512 3240 15564
rect 3292 15512 3298 15564
rect 8662 15552 8668 15564
rect 8220 15524 8668 15552
rect 2547 15456 2636 15484
rect 2685 15487 2743 15493
rect 2547 15453 2559 15456
rect 2501 15447 2559 15453
rect 2685 15453 2697 15487
rect 2731 15453 2743 15487
rect 2685 15447 2743 15453
rect 3050 15444 3056 15496
rect 3108 15484 3114 15496
rect 3145 15487 3203 15493
rect 3145 15484 3157 15487
rect 3108 15456 3157 15484
rect 3108 15444 3114 15456
rect 3145 15453 3157 15456
rect 3191 15453 3203 15487
rect 3145 15447 3203 15453
rect 3878 15444 3884 15496
rect 3936 15444 3942 15496
rect 6086 15444 6092 15496
rect 6144 15484 6150 15496
rect 6482 15487 6540 15493
rect 6482 15484 6494 15487
rect 6144 15456 6494 15484
rect 6144 15444 6150 15456
rect 6482 15453 6494 15456
rect 6528 15453 6540 15487
rect 6482 15447 6540 15453
rect 8018 15444 8024 15496
rect 8076 15444 8082 15496
rect 8220 15493 8248 15524
rect 8662 15512 8668 15524
rect 8720 15512 8726 15564
rect 9600 15561 9628 15592
rect 9766 15580 9772 15632
rect 9824 15620 9830 15632
rect 9953 15623 10011 15629
rect 9953 15620 9965 15623
rect 9824 15592 9965 15620
rect 9824 15580 9830 15592
rect 9953 15589 9965 15592
rect 9999 15620 10011 15623
rect 10410 15620 10416 15632
rect 9999 15592 10416 15620
rect 9999 15589 10011 15592
rect 9953 15583 10011 15589
rect 10410 15580 10416 15592
rect 10468 15580 10474 15632
rect 10520 15629 10548 15660
rect 11054 15648 11060 15700
rect 11112 15688 11118 15700
rect 11149 15691 11207 15697
rect 11149 15688 11161 15691
rect 11112 15660 11161 15688
rect 11112 15648 11118 15660
rect 11149 15657 11161 15660
rect 11195 15657 11207 15691
rect 11149 15651 11207 15657
rect 12713 15691 12771 15697
rect 12713 15657 12725 15691
rect 12759 15688 12771 15691
rect 12894 15688 12900 15700
rect 12759 15660 12900 15688
rect 12759 15657 12771 15660
rect 12713 15651 12771 15657
rect 12894 15648 12900 15660
rect 12952 15648 12958 15700
rect 10505 15623 10563 15629
rect 10505 15589 10517 15623
rect 10551 15620 10563 15623
rect 10962 15620 10968 15632
rect 10551 15592 10968 15620
rect 10551 15589 10563 15592
rect 10505 15583 10563 15589
rect 10962 15580 10968 15592
rect 11020 15580 11026 15632
rect 12434 15620 12440 15632
rect 11072 15592 12440 15620
rect 9585 15555 9643 15561
rect 9585 15521 9597 15555
rect 9631 15552 9643 15555
rect 9631 15524 10180 15552
rect 9631 15521 9643 15524
rect 9585 15515 9643 15521
rect 8205 15487 8263 15493
rect 8205 15453 8217 15487
rect 8251 15453 8263 15487
rect 8205 15447 8263 15453
rect 8481 15487 8539 15493
rect 8481 15453 8493 15487
rect 8527 15484 8539 15487
rect 8570 15484 8576 15496
rect 8527 15456 8576 15484
rect 8527 15453 8539 15456
rect 8481 15447 8539 15453
rect 8570 15444 8576 15456
rect 8628 15484 8634 15496
rect 9125 15487 9183 15493
rect 9125 15484 9137 15487
rect 8628 15456 9137 15484
rect 8628 15444 8634 15456
rect 9125 15453 9137 15456
rect 9171 15453 9183 15487
rect 9125 15447 9183 15453
rect 9398 15444 9404 15496
rect 9456 15484 9462 15496
rect 9769 15487 9827 15493
rect 9769 15484 9781 15487
rect 9456 15456 9781 15484
rect 9456 15444 9462 15456
rect 9769 15453 9781 15456
rect 9815 15453 9827 15487
rect 10152 15484 10180 15524
rect 10226 15512 10232 15564
rect 10284 15552 10290 15564
rect 10689 15555 10747 15561
rect 10689 15552 10701 15555
rect 10284 15524 10701 15552
rect 10284 15512 10290 15524
rect 10689 15521 10701 15524
rect 10735 15552 10747 15555
rect 11072 15552 11100 15592
rect 12434 15580 12440 15592
rect 12492 15580 12498 15632
rect 12805 15623 12863 15629
rect 12805 15589 12817 15623
rect 12851 15620 12863 15623
rect 13078 15620 13084 15632
rect 12851 15592 13084 15620
rect 12851 15589 12863 15592
rect 12805 15583 12863 15589
rect 13078 15580 13084 15592
rect 13136 15580 13142 15632
rect 13449 15623 13507 15629
rect 13449 15589 13461 15623
rect 13495 15589 13507 15623
rect 13449 15583 13507 15589
rect 10735 15524 11100 15552
rect 10735 15521 10747 15524
rect 10689 15515 10747 15521
rect 11072 15493 11100 15524
rect 11330 15512 11336 15564
rect 11388 15552 11394 15564
rect 11425 15555 11483 15561
rect 11425 15552 11437 15555
rect 11388 15524 11437 15552
rect 11388 15512 11394 15524
rect 11425 15521 11437 15524
rect 11471 15552 11483 15555
rect 13464 15552 13492 15583
rect 11471 15524 13492 15552
rect 11471 15521 11483 15524
rect 11425 15515 11483 15521
rect 13722 15512 13728 15564
rect 13780 15552 13786 15564
rect 14461 15555 14519 15561
rect 14461 15552 14473 15555
rect 13780 15524 14473 15552
rect 13780 15512 13786 15524
rect 14461 15521 14473 15524
rect 14507 15521 14519 15555
rect 14461 15515 14519 15521
rect 14550 15512 14556 15564
rect 14608 15552 14614 15564
rect 15565 15555 15623 15561
rect 15565 15552 15577 15555
rect 14608 15524 15577 15552
rect 14608 15512 14614 15524
rect 15565 15521 15577 15524
rect 15611 15521 15623 15555
rect 15565 15515 15623 15521
rect 16206 15512 16212 15564
rect 16264 15512 16270 15564
rect 11057 15487 11115 15493
rect 10152 15456 11008 15484
rect 9769 15447 9827 15453
rect 4157 15419 4215 15425
rect 4157 15385 4169 15419
rect 4203 15385 4215 15419
rect 4157 15379 4215 15385
rect 2593 15351 2651 15357
rect 2593 15317 2605 15351
rect 2639 15348 2651 15351
rect 2958 15348 2964 15360
rect 2639 15320 2964 15348
rect 2639 15317 2651 15320
rect 2593 15311 2651 15317
rect 2958 15308 2964 15320
rect 3016 15308 3022 15360
rect 3513 15351 3571 15357
rect 3513 15317 3525 15351
rect 3559 15348 3571 15351
rect 4172 15348 4200 15379
rect 4614 15376 4620 15428
rect 4672 15376 4678 15428
rect 7193 15419 7251 15425
rect 7193 15385 7205 15419
rect 7239 15416 7251 15419
rect 8294 15416 8300 15428
rect 7239 15388 8300 15416
rect 7239 15385 7251 15388
rect 7193 15379 7251 15385
rect 8294 15376 8300 15388
rect 8352 15416 8358 15428
rect 8846 15416 8852 15428
rect 8352 15388 8852 15416
rect 8352 15376 8358 15388
rect 8846 15376 8852 15388
rect 8904 15376 8910 15428
rect 9309 15419 9367 15425
rect 9309 15385 9321 15419
rect 9355 15416 9367 15419
rect 9582 15416 9588 15428
rect 9355 15388 9588 15416
rect 9355 15385 9367 15388
rect 9309 15379 9367 15385
rect 9582 15376 9588 15388
rect 9640 15376 9646 15428
rect 3559 15320 4200 15348
rect 3559 15317 3571 15320
rect 3513 15311 3571 15317
rect 4982 15308 4988 15360
rect 5040 15348 5046 15360
rect 5629 15351 5687 15357
rect 5629 15348 5641 15351
rect 5040 15320 5641 15348
rect 5040 15308 5046 15320
rect 5629 15317 5641 15320
rect 5675 15317 5687 15351
rect 5629 15311 5687 15317
rect 8110 15308 8116 15360
rect 8168 15308 8174 15360
rect 9784 15348 9812 15447
rect 10229 15419 10287 15425
rect 10229 15385 10241 15419
rect 10275 15416 10287 15419
rect 10318 15416 10324 15428
rect 10275 15388 10324 15416
rect 10275 15385 10287 15388
rect 10229 15379 10287 15385
rect 10318 15376 10324 15388
rect 10376 15376 10382 15428
rect 10980 15416 11008 15456
rect 11057 15453 11069 15487
rect 11103 15453 11115 15487
rect 11238 15484 11244 15496
rect 11057 15447 11115 15453
rect 11164 15456 11244 15484
rect 11164 15416 11192 15456
rect 11238 15444 11244 15456
rect 11296 15444 11302 15496
rect 11698 15444 11704 15496
rect 11756 15444 11762 15496
rect 11882 15444 11888 15496
rect 11940 15444 11946 15496
rect 12253 15487 12311 15493
rect 12253 15453 12265 15487
rect 12299 15453 12311 15487
rect 12253 15447 12311 15453
rect 12345 15487 12403 15493
rect 12345 15453 12357 15487
rect 12391 15484 12403 15487
rect 12710 15484 12716 15496
rect 12391 15456 12716 15484
rect 12391 15453 12403 15456
rect 12345 15447 12403 15453
rect 12268 15416 12296 15447
rect 12710 15444 12716 15456
rect 12768 15444 12774 15496
rect 13630 15444 13636 15496
rect 13688 15484 13694 15496
rect 14185 15487 14243 15493
rect 14185 15484 14197 15487
rect 13688 15456 14197 15484
rect 13688 15444 13694 15456
rect 14185 15453 14197 15456
rect 14231 15453 14243 15487
rect 14185 15447 14243 15453
rect 16485 15487 16543 15493
rect 16485 15453 16497 15487
rect 16531 15484 16543 15487
rect 16574 15484 16580 15496
rect 16531 15456 16580 15484
rect 16531 15453 16543 15456
rect 16485 15447 16543 15453
rect 16574 15444 16580 15456
rect 16632 15444 16638 15496
rect 13078 15416 13084 15428
rect 10980 15388 11192 15416
rect 11256 15388 11652 15416
rect 12268 15388 13084 15416
rect 10134 15348 10140 15360
rect 9784 15320 10140 15348
rect 10134 15308 10140 15320
rect 10192 15348 10198 15360
rect 11146 15348 11152 15360
rect 10192 15320 11152 15348
rect 10192 15308 10198 15320
rect 11146 15308 11152 15320
rect 11204 15308 11210 15360
rect 11256 15357 11284 15388
rect 11241 15351 11299 15357
rect 11241 15317 11253 15351
rect 11287 15317 11299 15351
rect 11624 15348 11652 15388
rect 13078 15376 13084 15388
rect 13136 15376 13142 15428
rect 13170 15376 13176 15428
rect 13228 15376 13234 15428
rect 12802 15348 12808 15360
rect 11624 15320 12808 15348
rect 11241 15311 11299 15317
rect 12802 15308 12808 15320
rect 12860 15308 12866 15360
rect 1104 15258 25852 15280
rect 1104 15206 8214 15258
rect 8266 15206 8278 15258
rect 8330 15206 8342 15258
rect 8394 15206 8406 15258
rect 8458 15206 8470 15258
rect 8522 15206 16214 15258
rect 16266 15206 16278 15258
rect 16330 15206 16342 15258
rect 16394 15206 16406 15258
rect 16458 15206 16470 15258
rect 16522 15206 24214 15258
rect 24266 15206 24278 15258
rect 24330 15206 24342 15258
rect 24394 15206 24406 15258
rect 24458 15206 24470 15258
rect 24522 15206 25852 15258
rect 1104 15184 25852 15206
rect 3878 15144 3884 15156
rect 1688 15116 3884 15144
rect 1486 14900 1492 14952
rect 1544 14940 1550 14952
rect 1688 14949 1716 15116
rect 3878 15104 3884 15116
rect 3936 15144 3942 15156
rect 6822 15144 6828 15156
rect 3936 15116 6828 15144
rect 3936 15104 3942 15116
rect 6822 15104 6828 15116
rect 6880 15104 6886 15156
rect 6932 15116 8432 15144
rect 2958 15036 2964 15088
rect 3016 15036 3022 15088
rect 3234 15036 3240 15088
rect 3292 15076 3298 15088
rect 4062 15076 4068 15088
rect 3292 15048 4068 15076
rect 3292 15036 3298 15048
rect 3712 15017 3740 15048
rect 4062 15036 4068 15048
rect 4120 15076 4126 15088
rect 6932 15076 6960 15116
rect 4120 15048 6960 15076
rect 4120 15036 4126 15048
rect 8110 15036 8116 15088
rect 8168 15036 8174 15088
rect 8404 15076 8432 15116
rect 8570 15104 8576 15156
rect 8628 15104 8634 15156
rect 10042 15104 10048 15156
rect 10100 15104 10106 15156
rect 10870 15104 10876 15156
rect 10928 15144 10934 15156
rect 11149 15147 11207 15153
rect 11149 15144 11161 15147
rect 10928 15116 11161 15144
rect 10928 15104 10934 15116
rect 11149 15113 11161 15116
rect 11195 15113 11207 15147
rect 11149 15107 11207 15113
rect 11422 15104 11428 15156
rect 11480 15144 11486 15156
rect 11609 15147 11667 15153
rect 11609 15144 11621 15147
rect 11480 15116 11621 15144
rect 11480 15104 11486 15116
rect 11609 15113 11621 15116
rect 11655 15113 11667 15147
rect 11609 15107 11667 15113
rect 11974 15104 11980 15156
rect 12032 15144 12038 15156
rect 12345 15147 12403 15153
rect 12345 15144 12357 15147
rect 12032 15116 12357 15144
rect 12032 15104 12038 15116
rect 12345 15113 12357 15116
rect 12391 15113 12403 15147
rect 12345 15107 12403 15113
rect 12802 15104 12808 15156
rect 12860 15104 12866 15156
rect 9858 15076 9864 15088
rect 8404 15048 9864 15076
rect 9858 15036 9864 15048
rect 9916 15036 9922 15088
rect 3697 15011 3755 15017
rect 3697 14977 3709 15011
rect 3743 14977 3755 15011
rect 3697 14971 3755 14977
rect 3881 15011 3939 15017
rect 3881 14977 3893 15011
rect 3927 15008 3939 15011
rect 3970 15008 3976 15020
rect 3927 14980 3976 15008
rect 3927 14977 3939 14980
rect 3881 14971 3939 14977
rect 3970 14968 3976 14980
rect 4028 14968 4034 15020
rect 4341 15011 4399 15017
rect 4341 14977 4353 15011
rect 4387 15008 4399 15011
rect 4798 15008 4804 15020
rect 4387 14980 4804 15008
rect 4387 14977 4399 14980
rect 4341 14971 4399 14977
rect 4798 14968 4804 14980
rect 4856 14968 4862 15020
rect 5353 15011 5411 15017
rect 5353 14977 5365 15011
rect 5399 14977 5411 15011
rect 5353 14971 5411 14977
rect 1673 14943 1731 14949
rect 1673 14940 1685 14943
rect 1544 14912 1685 14940
rect 1544 14900 1550 14912
rect 1673 14909 1685 14912
rect 1719 14909 1731 14943
rect 1673 14903 1731 14909
rect 1949 14943 2007 14949
rect 1949 14909 1961 14943
rect 1995 14940 2007 14943
rect 2682 14940 2688 14952
rect 1995 14912 2688 14940
rect 1995 14909 2007 14912
rect 1949 14903 2007 14909
rect 2682 14900 2688 14912
rect 2740 14900 2746 14952
rect 3234 14900 3240 14952
rect 3292 14940 3298 14952
rect 3789 14943 3847 14949
rect 3789 14940 3801 14943
rect 3292 14912 3801 14940
rect 3292 14900 3298 14912
rect 3789 14909 3801 14912
rect 3835 14909 3847 14943
rect 3789 14903 3847 14909
rect 4525 14943 4583 14949
rect 4525 14909 4537 14943
rect 4571 14940 4583 14943
rect 5074 14940 5080 14952
rect 4571 14912 5080 14940
rect 4571 14909 4583 14912
rect 4525 14903 4583 14909
rect 4540 14872 4568 14903
rect 5074 14900 5080 14912
rect 5132 14900 5138 14952
rect 5368 14940 5396 14971
rect 9122 14968 9128 15020
rect 9180 15008 9186 15020
rect 9493 15011 9551 15017
rect 9493 15008 9505 15011
rect 9180 14980 9505 15008
rect 9180 14968 9186 14980
rect 9493 14977 9505 14980
rect 9539 14977 9551 15011
rect 9493 14971 9551 14977
rect 10042 14968 10048 15020
rect 10100 14968 10106 15020
rect 10226 14968 10232 15020
rect 10284 14968 10290 15020
rect 11057 15011 11115 15017
rect 11057 14977 11069 15011
rect 11103 15008 11115 15011
rect 11146 15008 11152 15020
rect 11103 14980 11152 15008
rect 11103 14977 11115 14980
rect 11057 14971 11115 14977
rect 11146 14968 11152 14980
rect 11204 14968 11210 15020
rect 11238 14968 11244 15020
rect 11296 14968 11302 15020
rect 11330 14968 11336 15020
rect 11388 15008 11394 15020
rect 11609 15011 11667 15017
rect 11609 15008 11621 15011
rect 11388 14980 11621 15008
rect 11388 14968 11394 14980
rect 11609 14977 11621 14980
rect 11655 14977 11667 15011
rect 11609 14971 11667 14977
rect 11793 15011 11851 15017
rect 11793 14977 11805 15011
rect 11839 15008 11851 15011
rect 11992 15008 12020 15104
rect 13170 15076 13176 15088
rect 12452 15048 13176 15076
rect 11839 14980 12020 15008
rect 11839 14977 11851 14980
rect 11793 14971 11851 14977
rect 12066 14968 12072 15020
rect 12124 15008 12130 15020
rect 12452 15017 12480 15048
rect 13170 15036 13176 15048
rect 13228 15036 13234 15088
rect 16114 15036 16120 15088
rect 16172 15036 16178 15088
rect 12253 15011 12311 15017
rect 12253 15008 12265 15011
rect 12124 14980 12265 15008
rect 12124 14968 12130 14980
rect 12253 14977 12265 14980
rect 12299 14977 12311 15011
rect 12253 14971 12311 14977
rect 12437 15011 12495 15017
rect 12437 14977 12449 15011
rect 12483 14977 12495 15011
rect 12437 14971 12495 14977
rect 12713 15011 12771 15017
rect 12713 14977 12725 15011
rect 12759 14977 12771 15011
rect 12713 14971 12771 14977
rect 5368 14912 6776 14940
rect 3436 14844 4568 14872
rect 3436 14816 3464 14844
rect 4982 14832 4988 14884
rect 5040 14872 5046 14884
rect 5261 14875 5319 14881
rect 5261 14872 5273 14875
rect 5040 14844 5273 14872
rect 5040 14832 5046 14844
rect 5261 14841 5273 14844
rect 5307 14841 5319 14875
rect 5261 14835 5319 14841
rect 3418 14764 3424 14816
rect 3476 14764 3482 14816
rect 3510 14764 3516 14816
rect 3568 14804 3574 14816
rect 4157 14807 4215 14813
rect 4157 14804 4169 14807
rect 3568 14776 4169 14804
rect 3568 14764 3574 14776
rect 4157 14773 4169 14776
rect 4203 14773 4215 14807
rect 4157 14767 4215 14773
rect 5353 14807 5411 14813
rect 5353 14773 5365 14807
rect 5399 14804 5411 14807
rect 5718 14804 5724 14816
rect 5399 14776 5724 14804
rect 5399 14773 5411 14776
rect 5353 14767 5411 14773
rect 5718 14764 5724 14776
rect 5776 14764 5782 14816
rect 6748 14804 6776 14912
rect 6822 14900 6828 14952
rect 6880 14900 6886 14952
rect 7098 14900 7104 14952
rect 7156 14900 7162 14952
rect 9674 14900 9680 14952
rect 9732 14940 9738 14952
rect 9769 14943 9827 14949
rect 9769 14940 9781 14943
rect 9732 14912 9781 14940
rect 9732 14900 9738 14912
rect 9769 14909 9781 14912
rect 9815 14909 9827 14943
rect 11256 14940 11284 14968
rect 12728 14940 12756 14971
rect 13722 14968 13728 15020
rect 13780 14968 13786 15020
rect 16298 14968 16304 15020
rect 16356 14968 16362 15020
rect 16942 14968 16948 15020
rect 17000 14968 17006 15020
rect 11256 14912 12756 14940
rect 9769 14903 9827 14909
rect 15102 14900 15108 14952
rect 15160 14940 15166 14952
rect 15473 14943 15531 14949
rect 15473 14940 15485 14943
rect 15160 14912 15485 14940
rect 15160 14900 15166 14912
rect 15473 14909 15485 14912
rect 15519 14909 15531 14943
rect 15473 14903 15531 14909
rect 9306 14832 9312 14884
rect 9364 14872 9370 14884
rect 9364 14844 12434 14872
rect 9364 14832 9370 14844
rect 7834 14804 7840 14816
rect 6748 14776 7840 14804
rect 7834 14764 7840 14776
rect 7892 14764 7898 14816
rect 12406 14804 12434 14844
rect 12710 14832 12716 14884
rect 12768 14872 12774 14884
rect 13541 14875 13599 14881
rect 13541 14872 13553 14875
rect 12768 14844 13553 14872
rect 12768 14832 12774 14844
rect 13541 14841 13553 14844
rect 13587 14872 13599 14875
rect 13630 14872 13636 14884
rect 13587 14844 13636 14872
rect 13587 14841 13599 14844
rect 13541 14835 13599 14841
rect 13630 14832 13636 14844
rect 13688 14832 13694 14884
rect 12618 14804 12624 14816
rect 12406 14776 12624 14804
rect 12618 14764 12624 14776
rect 12676 14764 12682 14816
rect 16850 14764 16856 14816
rect 16908 14764 16914 14816
rect 1104 14714 25852 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 12214 14714
rect 12266 14662 12278 14714
rect 12330 14662 12342 14714
rect 12394 14662 12406 14714
rect 12458 14662 12470 14714
rect 12522 14662 20214 14714
rect 20266 14662 20278 14714
rect 20330 14662 20342 14714
rect 20394 14662 20406 14714
rect 20458 14662 20470 14714
rect 20522 14662 25852 14714
rect 1104 14640 25852 14662
rect 4062 14560 4068 14612
rect 4120 14600 4126 14612
rect 4120 14572 4384 14600
rect 4120 14560 4126 14572
rect 3050 14492 3056 14544
rect 3108 14532 3114 14544
rect 3108 14504 4200 14532
rect 3108 14492 3114 14504
rect 2130 14424 2136 14476
rect 2188 14464 2194 14476
rect 2188 14436 4108 14464
rect 2188 14424 2194 14436
rect 4080 14408 4108 14436
rect 1486 14356 1492 14408
rect 1544 14396 1550 14408
rect 1765 14399 1823 14405
rect 1765 14396 1777 14399
rect 1544 14368 1777 14396
rect 1544 14356 1550 14368
rect 1765 14365 1777 14368
rect 1811 14365 1823 14399
rect 1765 14359 1823 14365
rect 3142 14356 3148 14408
rect 3200 14356 3206 14408
rect 4062 14356 4068 14408
rect 4120 14356 4126 14408
rect 4172 14405 4200 14504
rect 4356 14405 4384 14572
rect 5074 14560 5080 14612
rect 5132 14560 5138 14612
rect 6825 14603 6883 14609
rect 6825 14569 6837 14603
rect 6871 14600 6883 14603
rect 7098 14600 7104 14612
rect 6871 14572 7104 14600
rect 6871 14569 6883 14572
rect 6825 14563 6883 14569
rect 7098 14560 7104 14572
rect 7156 14560 7162 14612
rect 8297 14603 8355 14609
rect 8297 14569 8309 14603
rect 8343 14600 8355 14603
rect 8662 14600 8668 14612
rect 8343 14572 8668 14600
rect 8343 14569 8355 14572
rect 8297 14563 8355 14569
rect 8662 14560 8668 14572
rect 8720 14600 8726 14612
rect 9674 14600 9680 14612
rect 8720 14572 9680 14600
rect 8720 14560 8726 14572
rect 9674 14560 9680 14572
rect 9732 14560 9738 14612
rect 9858 14560 9864 14612
rect 9916 14600 9922 14612
rect 9916 14572 12434 14600
rect 9916 14560 9922 14572
rect 5261 14535 5319 14541
rect 5261 14501 5273 14535
rect 5307 14532 5319 14535
rect 5307 14504 9720 14532
rect 5307 14501 5319 14504
rect 5261 14495 5319 14501
rect 6181 14467 6239 14473
rect 6181 14464 6193 14467
rect 4448 14436 6193 14464
rect 4448 14405 4476 14436
rect 6181 14433 6193 14436
rect 6227 14433 6239 14467
rect 8570 14464 8576 14476
rect 6181 14427 6239 14433
rect 7116 14436 8576 14464
rect 4157 14399 4215 14405
rect 4157 14365 4169 14399
rect 4203 14396 4215 14399
rect 4341 14399 4399 14405
rect 4203 14368 4292 14396
rect 4203 14365 4215 14368
rect 4157 14359 4215 14365
rect 2041 14331 2099 14337
rect 2041 14297 2053 14331
rect 2087 14297 2099 14331
rect 2041 14291 2099 14297
rect 2056 14260 2084 14291
rect 2958 14260 2964 14272
rect 2056 14232 2964 14260
rect 2958 14220 2964 14232
rect 3016 14220 3022 14272
rect 3513 14263 3571 14269
rect 3513 14229 3525 14263
rect 3559 14260 3571 14263
rect 3602 14260 3608 14272
rect 3559 14232 3608 14260
rect 3559 14229 3571 14232
rect 3513 14223 3571 14229
rect 3602 14220 3608 14232
rect 3660 14220 3666 14272
rect 3878 14220 3884 14272
rect 3936 14220 3942 14272
rect 4264 14260 4292 14368
rect 4341 14365 4353 14399
rect 4387 14365 4399 14399
rect 4341 14359 4399 14365
rect 4433 14399 4491 14405
rect 4433 14365 4445 14399
rect 4479 14365 4491 14399
rect 4433 14359 4491 14365
rect 4982 14356 4988 14408
rect 5040 14396 5046 14408
rect 5040 14368 6040 14396
rect 5040 14356 5046 14368
rect 4893 14331 4951 14337
rect 4893 14297 4905 14331
rect 4939 14328 4951 14331
rect 5258 14328 5264 14340
rect 4939 14300 5264 14328
rect 4939 14297 4951 14300
rect 4893 14291 4951 14297
rect 5258 14288 5264 14300
rect 5316 14288 5322 14340
rect 5350 14288 5356 14340
rect 5408 14328 5414 14340
rect 5629 14331 5687 14337
rect 5629 14328 5641 14331
rect 5408 14300 5641 14328
rect 5408 14288 5414 14300
rect 5629 14297 5641 14300
rect 5675 14297 5687 14331
rect 6012 14328 6040 14368
rect 6086 14356 6092 14408
rect 6144 14356 6150 14408
rect 6273 14399 6331 14405
rect 6273 14365 6285 14399
rect 6319 14365 6331 14399
rect 6273 14359 6331 14365
rect 6288 14328 6316 14359
rect 6638 14356 6644 14408
rect 6696 14356 6702 14408
rect 7116 14405 7144 14436
rect 8570 14424 8576 14436
rect 8628 14424 8634 14476
rect 9306 14424 9312 14476
rect 9364 14424 9370 14476
rect 9692 14473 9720 14504
rect 11054 14492 11060 14544
rect 11112 14532 11118 14544
rect 11882 14532 11888 14544
rect 11112 14504 11888 14532
rect 11112 14492 11118 14504
rect 9677 14467 9735 14473
rect 9677 14433 9689 14467
rect 9723 14433 9735 14467
rect 9677 14427 9735 14433
rect 9766 14424 9772 14476
rect 9824 14424 9830 14476
rect 10778 14464 10784 14476
rect 10520 14436 10784 14464
rect 7101 14399 7159 14405
rect 7101 14365 7113 14399
rect 7147 14365 7159 14399
rect 7101 14359 7159 14365
rect 7282 14356 7288 14408
rect 7340 14356 7346 14408
rect 7561 14399 7619 14405
rect 7561 14365 7573 14399
rect 7607 14365 7619 14399
rect 7561 14359 7619 14365
rect 8481 14399 8539 14405
rect 8481 14365 8493 14399
rect 8527 14396 8539 14399
rect 8846 14396 8852 14408
rect 8527 14368 8852 14396
rect 8527 14365 8539 14368
rect 8481 14359 8539 14365
rect 6012 14300 6316 14328
rect 5629 14291 5687 14297
rect 6822 14288 6828 14340
rect 6880 14328 6886 14340
rect 7576 14328 7604 14359
rect 8846 14356 8852 14368
rect 8904 14356 8910 14408
rect 9214 14356 9220 14408
rect 9272 14396 9278 14408
rect 9401 14399 9459 14405
rect 9401 14396 9413 14399
rect 9272 14368 9413 14396
rect 9272 14356 9278 14368
rect 9401 14365 9413 14368
rect 9447 14365 9459 14399
rect 9401 14359 9459 14365
rect 9539 14399 9597 14405
rect 9539 14365 9551 14399
rect 9585 14396 9597 14399
rect 10318 14396 10324 14408
rect 9585 14368 10324 14396
rect 9585 14365 9597 14368
rect 9539 14359 9597 14365
rect 10318 14356 10324 14368
rect 10376 14396 10382 14408
rect 10520 14405 10548 14436
rect 10778 14424 10784 14436
rect 10836 14424 10842 14476
rect 11517 14467 11575 14473
rect 11517 14464 11529 14467
rect 10980 14436 11529 14464
rect 10980 14405 11008 14436
rect 11517 14433 11529 14436
rect 11563 14433 11575 14467
rect 11517 14427 11575 14433
rect 11624 14405 11652 14504
rect 11882 14492 11888 14504
rect 11940 14492 11946 14544
rect 12406 14532 12434 14572
rect 12618 14560 12624 14612
rect 12676 14600 12682 14612
rect 13722 14600 13728 14612
rect 12676 14572 13728 14600
rect 12676 14560 12682 14572
rect 13722 14560 13728 14572
rect 13780 14600 13786 14612
rect 14645 14603 14703 14609
rect 14645 14600 14657 14603
rect 13780 14572 14657 14600
rect 13780 14560 13786 14572
rect 14645 14569 14657 14572
rect 14691 14569 14703 14603
rect 14645 14563 14703 14569
rect 15657 14603 15715 14609
rect 15657 14569 15669 14603
rect 15703 14600 15715 14603
rect 15746 14600 15752 14612
rect 15703 14572 15752 14600
rect 15703 14569 15715 14572
rect 15657 14563 15715 14569
rect 15746 14560 15752 14572
rect 15804 14560 15810 14612
rect 16853 14603 16911 14609
rect 16853 14569 16865 14603
rect 16899 14600 16911 14603
rect 16942 14600 16948 14612
rect 16899 14572 16948 14600
rect 16899 14569 16911 14572
rect 16853 14563 16911 14569
rect 16942 14560 16948 14572
rect 17000 14560 17006 14612
rect 12805 14535 12863 14541
rect 12805 14532 12817 14535
rect 12406 14504 12817 14532
rect 12805 14501 12817 14504
rect 12851 14501 12863 14535
rect 12805 14495 12863 14501
rect 11900 14464 11928 14492
rect 13173 14467 13231 14473
rect 11900 14436 13032 14464
rect 10505 14399 10563 14405
rect 10505 14396 10517 14399
rect 10376 14368 10517 14396
rect 10376 14356 10382 14368
rect 10505 14365 10517 14368
rect 10551 14365 10563 14399
rect 10505 14359 10563 14365
rect 10689 14399 10747 14405
rect 10689 14365 10701 14399
rect 10735 14396 10747 14399
rect 10965 14399 11023 14405
rect 10965 14396 10977 14399
rect 10735 14368 10977 14396
rect 10735 14365 10747 14368
rect 10689 14359 10747 14365
rect 10965 14365 10977 14368
rect 11011 14365 11023 14399
rect 10965 14359 11023 14365
rect 11149 14399 11207 14405
rect 11149 14365 11161 14399
rect 11195 14365 11207 14399
rect 11149 14359 11207 14365
rect 11609 14399 11667 14405
rect 11609 14365 11621 14399
rect 11655 14365 11667 14399
rect 11609 14359 11667 14365
rect 8938 14328 8944 14340
rect 6880 14300 8944 14328
rect 6880 14288 6886 14300
rect 8938 14288 8944 14300
rect 8996 14288 9002 14340
rect 9030 14288 9036 14340
rect 9088 14328 9094 14340
rect 10704 14328 10732 14359
rect 9088 14300 10732 14328
rect 9088 14288 9094 14300
rect 10778 14288 10784 14340
rect 10836 14328 10842 14340
rect 11164 14328 11192 14359
rect 12710 14356 12716 14408
rect 12768 14356 12774 14408
rect 12802 14356 12808 14408
rect 12860 14356 12866 14408
rect 12894 14356 12900 14408
rect 12952 14356 12958 14408
rect 13004 14405 13032 14436
rect 13173 14433 13185 14467
rect 13219 14464 13231 14467
rect 14458 14464 14464 14476
rect 13219 14436 14464 14464
rect 13219 14433 13231 14436
rect 13173 14427 13231 14433
rect 14458 14424 14464 14436
rect 14516 14424 14522 14476
rect 16298 14424 16304 14476
rect 16356 14424 16362 14476
rect 12989 14399 13047 14405
rect 12989 14365 13001 14399
rect 13035 14396 13047 14399
rect 13262 14396 13268 14408
rect 13035 14368 13268 14396
rect 13035 14365 13047 14368
rect 12989 14359 13047 14365
rect 13262 14356 13268 14368
rect 13320 14396 13326 14408
rect 13449 14399 13507 14405
rect 13449 14396 13461 14399
rect 13320 14368 13461 14396
rect 13320 14356 13326 14368
rect 13449 14365 13461 14368
rect 13495 14365 13507 14399
rect 13449 14359 13507 14365
rect 14182 14356 14188 14408
rect 14240 14356 14246 14408
rect 14829 14399 14887 14405
rect 14829 14365 14841 14399
rect 14875 14396 14887 14399
rect 15746 14396 15752 14408
rect 14875 14368 15752 14396
rect 14875 14365 14887 14368
rect 14829 14359 14887 14365
rect 15746 14356 15752 14368
rect 15804 14356 15810 14408
rect 15838 14356 15844 14408
rect 15896 14356 15902 14408
rect 16114 14356 16120 14408
rect 16172 14396 16178 14408
rect 16669 14399 16727 14405
rect 16669 14396 16681 14399
rect 16172 14368 16681 14396
rect 16172 14356 16178 14368
rect 16669 14365 16681 14368
rect 16715 14365 16727 14399
rect 16669 14359 16727 14365
rect 12618 14328 12624 14340
rect 10836 14300 12624 14328
rect 10836 14288 10842 14300
rect 12618 14288 12624 14300
rect 12676 14328 12682 14340
rect 13078 14328 13084 14340
rect 12676 14300 13084 14328
rect 12676 14288 12682 14300
rect 13078 14288 13084 14300
rect 13136 14288 13142 14340
rect 13170 14288 13176 14340
rect 13228 14328 13234 14340
rect 13633 14331 13691 14337
rect 13633 14328 13645 14331
rect 13228 14300 13645 14328
rect 13228 14288 13234 14300
rect 13633 14297 13645 14300
rect 13679 14328 13691 14331
rect 13679 14300 15700 14328
rect 13679 14297 13691 14300
rect 13633 14291 13691 14297
rect 4982 14260 4988 14272
rect 4264 14232 4988 14260
rect 4982 14220 4988 14232
rect 5040 14260 5046 14272
rect 5098 14263 5156 14269
rect 5098 14260 5110 14263
rect 5040 14232 5110 14260
rect 5040 14220 5046 14232
rect 5098 14229 5110 14232
rect 5144 14229 5156 14263
rect 5098 14223 5156 14229
rect 5721 14263 5779 14269
rect 5721 14229 5733 14263
rect 5767 14260 5779 14263
rect 5810 14260 5816 14272
rect 5767 14232 5816 14260
rect 5767 14229 5779 14232
rect 5721 14223 5779 14229
rect 5810 14220 5816 14232
rect 5868 14220 5874 14272
rect 7742 14220 7748 14272
rect 7800 14220 7806 14272
rect 9122 14220 9128 14272
rect 9180 14220 9186 14272
rect 10597 14263 10655 14269
rect 10597 14229 10609 14263
rect 10643 14260 10655 14263
rect 11054 14260 11060 14272
rect 10643 14232 11060 14260
rect 10643 14229 10655 14232
rect 10597 14223 10655 14229
rect 11054 14220 11060 14232
rect 11112 14220 11118 14272
rect 11149 14263 11207 14269
rect 11149 14229 11161 14263
rect 11195 14260 11207 14263
rect 11238 14260 11244 14272
rect 11195 14232 11244 14260
rect 11195 14229 11207 14232
rect 11149 14223 11207 14229
rect 11238 14220 11244 14232
rect 11296 14220 11302 14272
rect 11974 14220 11980 14272
rect 12032 14220 12038 14272
rect 14366 14220 14372 14272
rect 14424 14220 14430 14272
rect 15672 14269 15700 14300
rect 15657 14263 15715 14269
rect 15657 14229 15669 14263
rect 15703 14229 15715 14263
rect 15657 14223 15715 14229
rect 1104 14170 25852 14192
rect 1104 14118 8214 14170
rect 8266 14118 8278 14170
rect 8330 14118 8342 14170
rect 8394 14118 8406 14170
rect 8458 14118 8470 14170
rect 8522 14118 16214 14170
rect 16266 14118 16278 14170
rect 16330 14118 16342 14170
rect 16394 14118 16406 14170
rect 16458 14118 16470 14170
rect 16522 14118 24214 14170
rect 24266 14118 24278 14170
rect 24330 14118 24342 14170
rect 24394 14118 24406 14170
rect 24458 14118 24470 14170
rect 24522 14118 25852 14170
rect 1104 14096 25852 14118
rect 2225 14059 2283 14065
rect 2225 14025 2237 14059
rect 2271 14056 2283 14059
rect 3050 14056 3056 14068
rect 2271 14028 3056 14056
rect 2271 14025 2283 14028
rect 2225 14019 2283 14025
rect 3050 14016 3056 14028
rect 3108 14016 3114 14068
rect 3329 14059 3387 14065
rect 3329 14025 3341 14059
rect 3375 14056 3387 14059
rect 3878 14056 3884 14068
rect 3375 14028 3884 14056
rect 3375 14025 3387 14028
rect 3329 14019 3387 14025
rect 3878 14016 3884 14028
rect 3936 14016 3942 14068
rect 5258 14056 5264 14068
rect 3987 14028 5264 14056
rect 2409 13991 2467 13997
rect 2409 13957 2421 13991
rect 2455 13988 2467 13991
rect 3510 13988 3516 14000
rect 2455 13960 3516 13988
rect 2455 13957 2467 13960
rect 2409 13951 2467 13957
rect 3510 13948 3516 13960
rect 3568 13948 3574 14000
rect 3602 13948 3608 14000
rect 3660 13988 3666 14000
rect 3987 13988 4015 14028
rect 5258 14016 5264 14028
rect 5316 14016 5322 14068
rect 6638 14016 6644 14068
rect 6696 14056 6702 14068
rect 7101 14059 7159 14065
rect 7101 14056 7113 14059
rect 6696 14028 7113 14056
rect 6696 14016 6702 14028
rect 7101 14025 7113 14028
rect 7147 14025 7159 14059
rect 7101 14019 7159 14025
rect 7742 14016 7748 14068
rect 7800 14056 7806 14068
rect 16850 14056 16856 14068
rect 7800 14028 10364 14056
rect 7800 14016 7806 14028
rect 3660 13960 4015 13988
rect 3660 13948 3666 13960
rect 4062 13948 4068 14000
rect 4120 13988 4126 14000
rect 6086 13988 6092 14000
rect 4120 13960 6092 13988
rect 4120 13948 4126 13960
rect 2130 13880 2136 13932
rect 2188 13880 2194 13932
rect 4154 13920 4160 13932
rect 2424 13892 4160 13920
rect 2424 13793 2452 13892
rect 4154 13880 4160 13892
rect 4212 13920 4218 13932
rect 4249 13923 4307 13929
rect 4249 13920 4261 13923
rect 4212 13892 4261 13920
rect 4212 13880 4218 13892
rect 4249 13889 4261 13892
rect 4295 13889 4307 13923
rect 4893 13923 4951 13929
rect 4893 13920 4905 13923
rect 4249 13883 4307 13889
rect 4724 13892 4905 13920
rect 2682 13812 2688 13864
rect 2740 13812 2746 13864
rect 2869 13855 2927 13861
rect 2869 13821 2881 13855
rect 2915 13821 2927 13855
rect 2869 13815 2927 13821
rect 2961 13855 3019 13861
rect 2961 13821 2973 13855
rect 3007 13852 3019 13855
rect 3418 13852 3424 13864
rect 3007 13824 3424 13852
rect 3007 13821 3019 13824
rect 2961 13815 3019 13821
rect 2409 13787 2467 13793
rect 2409 13753 2421 13787
rect 2455 13753 2467 13787
rect 2884 13784 2912 13815
rect 3418 13812 3424 13824
rect 3476 13852 3482 13864
rect 4341 13855 4399 13861
rect 3476 13824 4292 13852
rect 3476 13812 3482 13824
rect 3326 13784 3332 13796
rect 2884 13756 3332 13784
rect 2409 13747 2467 13753
rect 3326 13744 3332 13756
rect 3384 13744 3390 13796
rect 4264 13784 4292 13824
rect 4341 13821 4353 13855
rect 4387 13852 4399 13855
rect 4614 13852 4620 13864
rect 4387 13824 4620 13852
rect 4387 13821 4399 13824
rect 4341 13815 4399 13821
rect 4614 13812 4620 13824
rect 4672 13812 4678 13864
rect 4724 13784 4752 13892
rect 4893 13889 4905 13892
rect 4939 13889 4951 13923
rect 4893 13883 4951 13889
rect 4798 13812 4804 13864
rect 4856 13812 4862 13864
rect 5092 13852 5120 13960
rect 6086 13948 6092 13960
rect 6144 13948 6150 14000
rect 6822 13948 6828 14000
rect 6880 13948 6886 14000
rect 8294 13988 8300 14000
rect 7392 13960 8300 13988
rect 5258 13880 5264 13932
rect 5316 13920 5322 13932
rect 5629 13923 5687 13929
rect 5629 13920 5641 13923
rect 5316 13892 5641 13920
rect 5316 13880 5322 13892
rect 5629 13889 5641 13892
rect 5675 13889 5687 13923
rect 5629 13883 5687 13889
rect 5718 13880 5724 13932
rect 5776 13880 5782 13932
rect 5810 13880 5816 13932
rect 5868 13920 5874 13932
rect 6641 13923 6699 13929
rect 6641 13920 6653 13923
rect 5868 13892 6653 13920
rect 5868 13880 5874 13892
rect 6641 13889 6653 13892
rect 6687 13920 6699 13923
rect 7392 13920 7420 13960
rect 8294 13948 8300 13960
rect 8352 13948 8358 14000
rect 9122 13988 9128 14000
rect 8404 13960 9128 13988
rect 6687 13892 7420 13920
rect 6687 13889 6699 13892
rect 6641 13883 6699 13889
rect 7466 13880 7472 13932
rect 7524 13880 7530 13932
rect 8404 13929 8432 13960
rect 9122 13948 9128 13960
rect 9180 13948 9186 14000
rect 9309 13991 9367 13997
rect 9309 13957 9321 13991
rect 9355 13988 9367 13991
rect 9858 13988 9864 14000
rect 9355 13960 9864 13988
rect 9355 13957 9367 13960
rect 9309 13951 9367 13957
rect 9858 13948 9864 13960
rect 9916 13948 9922 14000
rect 8388 13923 8446 13929
rect 8388 13889 8400 13923
rect 8434 13889 8446 13923
rect 8388 13883 8446 13889
rect 8478 13880 8484 13932
rect 8536 13880 8542 13932
rect 8570 13880 8576 13932
rect 8628 13920 8634 13932
rect 8757 13923 8815 13929
rect 8757 13920 8769 13923
rect 8628 13892 8769 13920
rect 8628 13880 8634 13892
rect 8757 13889 8769 13892
rect 8803 13889 8815 13923
rect 8757 13883 8815 13889
rect 8938 13880 8944 13932
rect 8996 13880 9002 13932
rect 9490 13880 9496 13932
rect 9548 13880 9554 13932
rect 10336 13929 10364 14028
rect 14108 14028 16856 14056
rect 11241 13991 11299 13997
rect 11241 13957 11253 13991
rect 11287 13988 11299 13991
rect 11287 13960 11928 13988
rect 11287 13957 11299 13960
rect 11241 13951 11299 13957
rect 10321 13923 10379 13929
rect 10321 13889 10333 13923
rect 10367 13889 10379 13923
rect 10321 13883 10379 13889
rect 10965 13923 11023 13929
rect 10965 13889 10977 13923
rect 11011 13920 11023 13923
rect 11054 13920 11060 13932
rect 11011 13892 11060 13920
rect 11011 13889 11023 13892
rect 10965 13883 11023 13889
rect 6457 13855 6515 13861
rect 5092 13824 5304 13852
rect 5276 13793 5304 13824
rect 6457 13821 6469 13855
rect 6503 13852 6515 13855
rect 7558 13852 7564 13864
rect 6503 13824 7564 13852
rect 6503 13821 6515 13824
rect 6457 13815 6515 13821
rect 7558 13812 7564 13824
rect 7616 13812 7622 13864
rect 7745 13855 7803 13861
rect 7745 13821 7757 13855
rect 7791 13852 7803 13855
rect 9508 13852 9536 13880
rect 7791 13824 9536 13852
rect 7791 13821 7803 13824
rect 7745 13815 7803 13821
rect 4264 13756 4752 13784
rect 5261 13787 5319 13793
rect 5261 13753 5273 13787
rect 5307 13753 5319 13787
rect 5261 13747 5319 13753
rect 7098 13744 7104 13796
rect 7156 13784 7162 13796
rect 8113 13787 8171 13793
rect 8113 13784 8125 13787
rect 7156 13756 8125 13784
rect 7156 13744 7162 13756
rect 8113 13753 8125 13756
rect 8159 13753 8171 13787
rect 8113 13747 8171 13753
rect 8478 13744 8484 13796
rect 8536 13784 8542 13796
rect 9030 13784 9036 13796
rect 8536 13756 9036 13784
rect 8536 13744 8542 13756
rect 9030 13744 9036 13756
rect 9088 13744 9094 13796
rect 10336 13784 10364 13883
rect 11054 13880 11060 13892
rect 11112 13880 11118 13932
rect 11900 13929 11928 13960
rect 14108 13932 14136 14028
rect 16850 14016 16856 14028
rect 16908 14016 16914 14068
rect 14366 13948 14372 14000
rect 14424 13948 14430 14000
rect 11885 13923 11943 13929
rect 11885 13889 11897 13923
rect 11931 13920 11943 13923
rect 12894 13920 12900 13932
rect 11931 13892 12900 13920
rect 11931 13889 11943 13892
rect 11885 13883 11943 13889
rect 12894 13880 12900 13892
rect 12952 13880 12958 13932
rect 14090 13880 14096 13932
rect 14148 13880 14154 13932
rect 15470 13880 15476 13932
rect 15528 13880 15534 13932
rect 16301 13923 16359 13929
rect 16301 13889 16313 13923
rect 16347 13920 16359 13923
rect 16758 13920 16764 13932
rect 16347 13892 16764 13920
rect 16347 13889 16359 13892
rect 16301 13883 16359 13889
rect 16758 13880 16764 13892
rect 16816 13880 16822 13932
rect 10413 13855 10471 13861
rect 10413 13821 10425 13855
rect 10459 13852 10471 13855
rect 11146 13852 11152 13864
rect 10459 13824 11152 13852
rect 10459 13821 10471 13824
rect 10413 13815 10471 13821
rect 11146 13812 11152 13824
rect 11204 13812 11210 13864
rect 11238 13812 11244 13864
rect 11296 13812 11302 13864
rect 11974 13812 11980 13864
rect 12032 13812 12038 13864
rect 12066 13812 12072 13864
rect 12124 13852 12130 13864
rect 12529 13855 12587 13861
rect 12529 13852 12541 13855
rect 12124 13824 12541 13852
rect 12124 13812 12130 13824
rect 12529 13821 12541 13824
rect 12575 13821 12587 13855
rect 12529 13815 12587 13821
rect 12618 13812 12624 13864
rect 12676 13852 12682 13864
rect 12805 13855 12863 13861
rect 12805 13852 12817 13855
rect 12676 13824 12817 13852
rect 12676 13812 12682 13824
rect 12805 13821 12817 13824
rect 12851 13821 12863 13855
rect 15102 13852 15108 13864
rect 12805 13815 12863 13821
rect 13740 13824 15108 13852
rect 11057 13787 11115 13793
rect 11057 13784 11069 13787
rect 10336 13756 11069 13784
rect 11057 13753 11069 13756
rect 11103 13753 11115 13787
rect 13740 13784 13768 13824
rect 15102 13812 15108 13824
rect 15160 13812 15166 13864
rect 15838 13812 15844 13864
rect 15896 13812 15902 13864
rect 11057 13747 11115 13753
rect 12084 13756 13768 13784
rect 3970 13676 3976 13728
rect 4028 13676 4034 13728
rect 5997 13719 6055 13725
rect 5997 13685 6009 13719
rect 6043 13716 6055 13719
rect 6454 13716 6460 13728
rect 6043 13688 6460 13716
rect 6043 13685 6055 13688
rect 5997 13679 6055 13685
rect 6454 13676 6460 13688
rect 6512 13676 6518 13728
rect 8754 13676 8760 13728
rect 8812 13676 8818 13728
rect 10502 13676 10508 13728
rect 10560 13716 10566 13728
rect 10597 13719 10655 13725
rect 10597 13716 10609 13719
rect 10560 13688 10609 13716
rect 10560 13676 10566 13688
rect 10597 13685 10609 13688
rect 10643 13685 10655 13719
rect 10597 13679 10655 13685
rect 10870 13676 10876 13728
rect 10928 13716 10934 13728
rect 12084 13716 12112 13756
rect 15378 13744 15384 13796
rect 15436 13784 15442 13796
rect 16117 13787 16175 13793
rect 16117 13784 16129 13787
rect 15436 13756 16129 13784
rect 15436 13744 15442 13756
rect 16117 13753 16129 13756
rect 16163 13753 16175 13787
rect 16117 13747 16175 13753
rect 10928 13688 12112 13716
rect 12161 13719 12219 13725
rect 10928 13676 10934 13688
rect 12161 13685 12173 13719
rect 12207 13716 12219 13719
rect 13354 13716 13360 13728
rect 12207 13688 13360 13716
rect 12207 13685 12219 13688
rect 12161 13679 12219 13685
rect 13354 13676 13360 13688
rect 13412 13676 13418 13728
rect 1104 13626 25852 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 12214 13626
rect 12266 13574 12278 13626
rect 12330 13574 12342 13626
rect 12394 13574 12406 13626
rect 12458 13574 12470 13626
rect 12522 13574 20214 13626
rect 20266 13574 20278 13626
rect 20330 13574 20342 13626
rect 20394 13574 20406 13626
rect 20458 13574 20470 13626
rect 20522 13574 25852 13626
rect 1104 13552 25852 13574
rect 2958 13472 2964 13524
rect 3016 13472 3022 13524
rect 7377 13515 7435 13521
rect 7377 13481 7389 13515
rect 7423 13512 7435 13515
rect 7466 13512 7472 13524
rect 7423 13484 7472 13512
rect 7423 13481 7435 13484
rect 7377 13475 7435 13481
rect 7466 13472 7472 13484
rect 7524 13472 7530 13524
rect 8297 13515 8355 13521
rect 8297 13481 8309 13515
rect 8343 13512 8355 13515
rect 8570 13512 8576 13524
rect 8343 13484 8576 13512
rect 8343 13481 8355 13484
rect 8297 13475 8355 13481
rect 8570 13472 8576 13484
rect 8628 13472 8634 13524
rect 11885 13515 11943 13521
rect 11885 13481 11897 13515
rect 11931 13512 11943 13515
rect 12066 13512 12072 13524
rect 11931 13484 12072 13512
rect 11931 13481 11943 13484
rect 11885 13475 11943 13481
rect 12066 13472 12072 13484
rect 12124 13472 12130 13524
rect 13725 13515 13783 13521
rect 13725 13481 13737 13515
rect 13771 13512 13783 13515
rect 14182 13512 14188 13524
rect 13771 13484 14188 13512
rect 13771 13481 13783 13484
rect 13725 13475 13783 13481
rect 14182 13472 14188 13484
rect 14240 13472 14246 13524
rect 15746 13472 15752 13524
rect 15804 13512 15810 13524
rect 15933 13515 15991 13521
rect 15933 13512 15945 13515
rect 15804 13484 15945 13512
rect 15804 13472 15810 13484
rect 15933 13481 15945 13484
rect 15979 13481 15991 13515
rect 15933 13475 15991 13481
rect 16022 13472 16028 13524
rect 16080 13512 16086 13524
rect 16761 13515 16819 13521
rect 16761 13512 16773 13515
rect 16080 13484 16773 13512
rect 16080 13472 16086 13484
rect 16761 13481 16773 13484
rect 16807 13481 16819 13515
rect 16761 13475 16819 13481
rect 4433 13447 4491 13453
rect 4433 13413 4445 13447
rect 4479 13444 4491 13447
rect 4614 13444 4620 13456
rect 4479 13416 4620 13444
rect 4479 13413 4491 13416
rect 4433 13407 4491 13413
rect 4614 13404 4620 13416
rect 4672 13404 4678 13456
rect 3326 13336 3332 13388
rect 3384 13376 3390 13388
rect 3384 13348 3464 13376
rect 3384 13336 3390 13348
rect 3145 13311 3203 13317
rect 3145 13277 3157 13311
rect 3191 13308 3203 13311
rect 3234 13308 3240 13320
rect 3191 13280 3240 13308
rect 3191 13277 3203 13280
rect 3145 13271 3203 13277
rect 3234 13268 3240 13280
rect 3292 13268 3298 13320
rect 3436 13317 3464 13348
rect 3878 13336 3884 13388
rect 3936 13376 3942 13388
rect 3973 13379 4031 13385
rect 3973 13376 3985 13379
rect 3936 13348 3985 13376
rect 3936 13336 3942 13348
rect 3973 13345 3985 13348
rect 4019 13376 4031 13379
rect 4798 13376 4804 13388
rect 4019 13348 4804 13376
rect 4019 13345 4031 13348
rect 3973 13339 4031 13345
rect 4798 13336 4804 13348
rect 4856 13376 4862 13388
rect 5077 13379 5135 13385
rect 4856 13348 4936 13376
rect 4856 13336 4862 13348
rect 3421 13311 3479 13317
rect 3421 13277 3433 13311
rect 3467 13277 3479 13311
rect 3421 13271 3479 13277
rect 3602 13268 3608 13320
rect 3660 13308 3666 13320
rect 4065 13311 4123 13317
rect 4065 13308 4077 13311
rect 3660 13280 4077 13308
rect 3660 13268 3666 13280
rect 4065 13277 4077 13280
rect 4111 13277 4123 13311
rect 4065 13271 4123 13277
rect 4706 13268 4712 13320
rect 4764 13268 4770 13320
rect 4908 13317 4936 13348
rect 5077 13345 5089 13379
rect 5123 13376 5135 13379
rect 5997 13379 6055 13385
rect 5123 13348 5856 13376
rect 5123 13345 5135 13348
rect 5077 13339 5135 13345
rect 4893 13311 4951 13317
rect 4893 13277 4905 13311
rect 4939 13308 4951 13311
rect 5258 13308 5264 13320
rect 4939 13280 5264 13308
rect 4939 13277 4951 13280
rect 4893 13271 4951 13277
rect 5258 13268 5264 13280
rect 5316 13268 5322 13320
rect 5350 13268 5356 13320
rect 5408 13268 5414 13320
rect 5534 13268 5540 13320
rect 5592 13268 5598 13320
rect 5828 13317 5856 13348
rect 5997 13345 6009 13379
rect 6043 13376 6055 13379
rect 7282 13376 7288 13388
rect 6043 13348 7288 13376
rect 6043 13345 6055 13348
rect 5997 13339 6055 13345
rect 7282 13336 7288 13348
rect 7340 13376 7346 13388
rect 7561 13379 7619 13385
rect 7561 13376 7573 13379
rect 7340 13348 7573 13376
rect 7340 13336 7346 13348
rect 7561 13345 7573 13348
rect 7607 13345 7619 13379
rect 8754 13376 8760 13388
rect 7561 13339 7619 13345
rect 7668 13348 8760 13376
rect 5813 13311 5871 13317
rect 5813 13277 5825 13311
rect 5859 13308 5871 13311
rect 6270 13308 6276 13320
rect 5859 13280 6276 13308
rect 5859 13277 5871 13280
rect 5813 13271 5871 13277
rect 6270 13268 6276 13280
rect 6328 13268 6334 13320
rect 6362 13268 6368 13320
rect 6420 13268 6426 13320
rect 6454 13268 6460 13320
rect 6512 13268 6518 13320
rect 6825 13311 6883 13317
rect 6825 13277 6837 13311
rect 6871 13308 6883 13311
rect 7098 13308 7104 13320
rect 6871 13280 7104 13308
rect 6871 13277 6883 13280
rect 6825 13271 6883 13277
rect 7098 13268 7104 13280
rect 7156 13268 7162 13320
rect 7668 13317 7696 13348
rect 8754 13336 8760 13348
rect 8812 13336 8818 13388
rect 10137 13379 10195 13385
rect 10137 13345 10149 13379
rect 10183 13376 10195 13379
rect 10410 13376 10416 13388
rect 10183 13348 10416 13376
rect 10183 13345 10195 13348
rect 10137 13339 10195 13345
rect 10410 13336 10416 13348
rect 10468 13336 10474 13388
rect 12802 13336 12808 13388
rect 12860 13376 12866 13388
rect 13081 13379 13139 13385
rect 13081 13376 13093 13379
rect 12860 13348 13093 13376
rect 12860 13336 12866 13348
rect 13081 13345 13093 13348
rect 13127 13345 13139 13379
rect 13081 13339 13139 13345
rect 13262 13336 13268 13388
rect 13320 13336 13326 13388
rect 14090 13336 14096 13388
rect 14148 13376 14154 13388
rect 14185 13379 14243 13385
rect 14185 13376 14197 13379
rect 14148 13348 14197 13376
rect 14148 13336 14154 13348
rect 14185 13345 14197 13348
rect 14231 13345 14243 13379
rect 14185 13339 14243 13345
rect 14458 13336 14464 13388
rect 14516 13336 14522 13388
rect 7653 13311 7711 13317
rect 7653 13277 7665 13311
rect 7699 13277 7711 13311
rect 7653 13271 7711 13277
rect 8113 13311 8171 13317
rect 8113 13277 8125 13311
rect 8159 13277 8171 13311
rect 8113 13271 8171 13277
rect 8297 13311 8355 13317
rect 8297 13277 8309 13311
rect 8343 13308 8355 13311
rect 8478 13308 8484 13320
rect 8343 13280 8484 13308
rect 8343 13277 8355 13280
rect 8297 13271 8355 13277
rect 3329 13243 3387 13249
rect 3329 13209 3341 13243
rect 3375 13240 3387 13243
rect 3620 13240 3648 13268
rect 3375 13212 3648 13240
rect 4724 13240 4752 13268
rect 6730 13240 6736 13252
rect 4724 13212 6736 13240
rect 3375 13209 3387 13212
rect 3329 13203 3387 13209
rect 6730 13200 6736 13212
rect 6788 13200 6794 13252
rect 7006 13200 7012 13252
rect 7064 13200 7070 13252
rect 7558 13200 7564 13252
rect 7616 13240 7622 13252
rect 8128 13240 8156 13271
rect 8478 13268 8484 13280
rect 8536 13268 8542 13320
rect 9214 13268 9220 13320
rect 9272 13268 9278 13320
rect 9582 13308 9588 13320
rect 9324 13280 9588 13308
rect 9324 13240 9352 13280
rect 9582 13268 9588 13280
rect 9640 13268 9646 13320
rect 9674 13268 9680 13320
rect 9732 13268 9738 13320
rect 9858 13268 9864 13320
rect 9916 13268 9922 13320
rect 13354 13268 13360 13320
rect 13412 13268 13418 13320
rect 16669 13311 16727 13317
rect 16669 13277 16681 13311
rect 16715 13308 16727 13311
rect 16758 13308 16764 13320
rect 16715 13280 16764 13308
rect 16715 13277 16727 13280
rect 16669 13271 16727 13277
rect 16758 13268 16764 13280
rect 16816 13268 16822 13320
rect 10413 13243 10471 13249
rect 10413 13240 10425 13243
rect 7616 13212 9352 13240
rect 9416 13212 10425 13240
rect 7616 13200 7622 13212
rect 9416 13181 9444 13212
rect 10413 13209 10425 13212
rect 10459 13209 10471 13243
rect 10413 13203 10471 13209
rect 10520 13212 10902 13240
rect 9401 13175 9459 13181
rect 9401 13141 9413 13175
rect 9447 13141 9459 13175
rect 9401 13135 9459 13141
rect 9769 13175 9827 13181
rect 9769 13141 9781 13175
rect 9815 13172 9827 13175
rect 10520 13172 10548 13212
rect 15010 13200 15016 13252
rect 15068 13200 15074 13252
rect 9815 13144 10548 13172
rect 9815 13141 9827 13144
rect 9769 13135 9827 13141
rect 1104 13082 25852 13104
rect 1104 13030 8214 13082
rect 8266 13030 8278 13082
rect 8330 13030 8342 13082
rect 8394 13030 8406 13082
rect 8458 13030 8470 13082
rect 8522 13030 16214 13082
rect 16266 13030 16278 13082
rect 16330 13030 16342 13082
rect 16394 13030 16406 13082
rect 16458 13030 16470 13082
rect 16522 13030 24214 13082
rect 24266 13030 24278 13082
rect 24330 13030 24342 13082
rect 24394 13030 24406 13082
rect 24458 13030 24470 13082
rect 24522 13030 25852 13082
rect 1104 13008 25852 13030
rect 6089 12971 6147 12977
rect 6089 12937 6101 12971
rect 6135 12968 6147 12971
rect 7469 12971 7527 12977
rect 7469 12968 7481 12971
rect 6135 12940 7481 12968
rect 6135 12937 6147 12940
rect 6089 12931 6147 12937
rect 7469 12937 7481 12940
rect 7515 12937 7527 12971
rect 7469 12931 7527 12937
rect 8846 12928 8852 12980
rect 8904 12928 8910 12980
rect 9214 12928 9220 12980
rect 9272 12968 9278 12980
rect 10137 12971 10195 12977
rect 10137 12968 10149 12971
rect 9272 12940 10149 12968
rect 9272 12928 9278 12940
rect 10137 12937 10149 12940
rect 10183 12937 10195 12971
rect 10137 12931 10195 12937
rect 10502 12928 10508 12980
rect 10560 12928 10566 12980
rect 10597 12971 10655 12977
rect 10597 12937 10609 12971
rect 10643 12968 10655 12971
rect 10778 12968 10784 12980
rect 10643 12940 10784 12968
rect 10643 12937 10655 12940
rect 10597 12931 10655 12937
rect 10778 12928 10784 12940
rect 10836 12928 10842 12980
rect 11146 12928 11152 12980
rect 11204 12968 11210 12980
rect 11609 12971 11667 12977
rect 11609 12968 11621 12971
rect 11204 12940 11621 12968
rect 11204 12928 11210 12940
rect 11609 12937 11621 12940
rect 11655 12937 11667 12971
rect 11609 12931 11667 12937
rect 15010 12928 15016 12980
rect 15068 12928 15074 12980
rect 15470 12928 15476 12980
rect 15528 12928 15534 12980
rect 3881 12903 3939 12909
rect 3881 12869 3893 12903
rect 3927 12900 3939 12903
rect 5169 12903 5227 12909
rect 3927 12872 4568 12900
rect 3927 12869 3939 12872
rect 3881 12863 3939 12869
rect 3602 12792 3608 12844
rect 3660 12832 3666 12844
rect 3789 12835 3847 12841
rect 3789 12832 3801 12835
rect 3660 12804 3801 12832
rect 3660 12792 3666 12804
rect 3789 12801 3801 12804
rect 3835 12801 3847 12835
rect 3973 12835 4031 12841
rect 3973 12832 3985 12835
rect 3789 12795 3847 12801
rect 3896 12804 3985 12832
rect 3896 12776 3924 12804
rect 3973 12801 3985 12804
rect 4019 12801 4031 12835
rect 3973 12795 4031 12801
rect 4154 12792 4160 12844
rect 4212 12832 4218 12844
rect 4540 12841 4568 12872
rect 5169 12869 5181 12903
rect 5215 12900 5227 12903
rect 5350 12900 5356 12912
rect 5215 12872 5356 12900
rect 5215 12869 5227 12872
rect 5169 12863 5227 12869
rect 5350 12860 5356 12872
rect 5408 12900 5414 12912
rect 5408 12872 6684 12900
rect 5408 12860 5414 12872
rect 4249 12835 4307 12841
rect 4249 12832 4261 12835
rect 4212 12804 4261 12832
rect 4212 12792 4218 12804
rect 4249 12801 4261 12804
rect 4295 12801 4307 12835
rect 4249 12795 4307 12801
rect 4525 12835 4583 12841
rect 4525 12801 4537 12835
rect 4571 12801 4583 12835
rect 4525 12795 4583 12801
rect 4706 12792 4712 12844
rect 4764 12832 4770 12844
rect 5077 12835 5135 12841
rect 5077 12832 5089 12835
rect 4764 12804 5089 12832
rect 4764 12792 4770 12804
rect 5077 12801 5089 12804
rect 5123 12801 5135 12835
rect 5077 12795 5135 12801
rect 5258 12792 5264 12844
rect 5316 12792 5322 12844
rect 5534 12792 5540 12844
rect 5592 12832 5598 12844
rect 5721 12835 5779 12841
rect 5721 12832 5733 12835
rect 5592 12804 5733 12832
rect 5592 12792 5598 12804
rect 5721 12801 5733 12804
rect 5767 12801 5779 12835
rect 5721 12795 5779 12801
rect 3878 12724 3884 12776
rect 3936 12724 3942 12776
rect 4341 12767 4399 12773
rect 4341 12733 4353 12767
rect 4387 12764 4399 12767
rect 4614 12764 4620 12776
rect 4387 12736 4620 12764
rect 4387 12733 4399 12736
rect 4341 12727 4399 12733
rect 4614 12724 4620 12736
rect 4672 12724 4678 12776
rect 4709 12631 4767 12637
rect 4709 12597 4721 12631
rect 4755 12628 4767 12631
rect 5736 12628 5764 12795
rect 6270 12792 6276 12844
rect 6328 12832 6334 12844
rect 6656 12841 6684 12872
rect 6730 12860 6736 12912
rect 6788 12900 6794 12912
rect 7377 12903 7435 12909
rect 7377 12900 7389 12903
rect 6788 12872 7389 12900
rect 6788 12860 6794 12872
rect 7377 12869 7389 12872
rect 7423 12900 7435 12903
rect 9398 12900 9404 12912
rect 7423 12872 9404 12900
rect 7423 12869 7435 12872
rect 7377 12863 7435 12869
rect 9398 12860 9404 12872
rect 9456 12900 9462 12912
rect 9585 12903 9643 12909
rect 9585 12900 9597 12903
rect 9456 12872 9597 12900
rect 9456 12860 9462 12872
rect 9585 12869 9597 12872
rect 9631 12869 9643 12903
rect 9585 12863 9643 12869
rect 9769 12903 9827 12909
rect 9769 12869 9781 12903
rect 9815 12900 9827 12903
rect 10042 12900 10048 12912
rect 9815 12872 10048 12900
rect 9815 12869 9827 12872
rect 9769 12863 9827 12869
rect 10042 12860 10048 12872
rect 10100 12860 10106 12912
rect 11054 12860 11060 12912
rect 11112 12900 11118 12912
rect 12069 12903 12127 12909
rect 12069 12900 12081 12903
rect 11112 12872 12081 12900
rect 11112 12860 11118 12872
rect 12069 12869 12081 12872
rect 12115 12869 12127 12903
rect 16022 12900 16028 12912
rect 12069 12863 12127 12869
rect 15120 12872 16028 12900
rect 6457 12835 6515 12841
rect 6457 12832 6469 12835
rect 6328 12804 6469 12832
rect 6328 12792 6334 12804
rect 6457 12801 6469 12804
rect 6503 12801 6515 12835
rect 6457 12795 6515 12801
rect 6641 12835 6699 12841
rect 6641 12801 6653 12835
rect 6687 12801 6699 12835
rect 8113 12835 8171 12841
rect 8113 12832 8125 12835
rect 6641 12795 6699 12801
rect 7852 12804 8125 12832
rect 5813 12767 5871 12773
rect 5813 12733 5825 12767
rect 5859 12764 5871 12767
rect 6549 12767 6607 12773
rect 6549 12764 6561 12767
rect 5859 12736 6561 12764
rect 5859 12733 5871 12736
rect 5813 12727 5871 12733
rect 6549 12733 6561 12736
rect 6595 12733 6607 12767
rect 6549 12727 6607 12733
rect 7006 12724 7012 12776
rect 7064 12764 7070 12776
rect 7285 12767 7343 12773
rect 7285 12764 7297 12767
rect 7064 12736 7297 12764
rect 7064 12724 7070 12736
rect 7285 12733 7297 12736
rect 7331 12733 7343 12767
rect 7285 12727 7343 12733
rect 7300 12696 7328 12727
rect 7852 12705 7880 12804
rect 8113 12801 8125 12804
rect 8159 12801 8171 12835
rect 8113 12795 8171 12801
rect 9033 12835 9091 12841
rect 9033 12801 9045 12835
rect 9079 12832 9091 12835
rect 9674 12832 9680 12844
rect 9079 12804 9680 12832
rect 9079 12801 9091 12804
rect 9033 12795 9091 12801
rect 9674 12792 9680 12804
rect 9732 12792 9738 12844
rect 9858 12792 9864 12844
rect 9916 12832 9922 12844
rect 10870 12832 10876 12844
rect 9916 12804 10876 12832
rect 9916 12792 9922 12804
rect 10870 12792 10876 12804
rect 10928 12792 10934 12844
rect 14921 12835 14979 12841
rect 14921 12801 14933 12835
rect 14967 12801 14979 12835
rect 14921 12795 14979 12801
rect 10689 12767 10747 12773
rect 10689 12733 10701 12767
rect 10735 12733 10747 12767
rect 10689 12727 10747 12733
rect 7837 12699 7895 12705
rect 7300 12668 7420 12696
rect 4755 12600 5764 12628
rect 7392 12628 7420 12668
rect 7837 12665 7849 12699
rect 7883 12665 7895 12699
rect 9490 12696 9496 12708
rect 7837 12659 7895 12665
rect 8128 12668 9496 12696
rect 8128 12628 8156 12668
rect 9490 12656 9496 12668
rect 9548 12696 9554 12708
rect 10704 12696 10732 12727
rect 14826 12724 14832 12776
rect 14884 12764 14890 12776
rect 14936 12764 14964 12795
rect 15010 12792 15016 12844
rect 15068 12832 15074 12844
rect 15120 12841 15148 12872
rect 15580 12841 15608 12872
rect 16022 12860 16028 12872
rect 16080 12900 16086 12912
rect 16080 12872 16988 12900
rect 16080 12860 16086 12872
rect 16960 12841 16988 12872
rect 15105 12835 15163 12841
rect 15105 12832 15117 12835
rect 15068 12804 15117 12832
rect 15068 12792 15074 12804
rect 15105 12801 15117 12804
rect 15151 12801 15163 12835
rect 15105 12795 15163 12801
rect 15381 12835 15439 12841
rect 15381 12801 15393 12835
rect 15427 12801 15439 12835
rect 15381 12795 15439 12801
rect 15565 12835 15623 12841
rect 15565 12801 15577 12835
rect 15611 12801 15623 12835
rect 15565 12795 15623 12801
rect 16761 12835 16819 12841
rect 16761 12801 16773 12835
rect 16807 12801 16819 12835
rect 16761 12795 16819 12801
rect 16945 12835 17003 12841
rect 16945 12801 16957 12835
rect 16991 12832 17003 12835
rect 17221 12835 17279 12841
rect 17221 12832 17233 12835
rect 16991 12804 17233 12832
rect 16991 12801 17003 12804
rect 16945 12795 17003 12801
rect 17221 12801 17233 12804
rect 17267 12801 17279 12835
rect 17221 12795 17279 12801
rect 17405 12835 17463 12841
rect 17405 12801 17417 12835
rect 17451 12832 17463 12835
rect 17862 12832 17868 12844
rect 17451 12804 17868 12832
rect 17451 12801 17463 12804
rect 17405 12795 17463 12801
rect 15396 12764 15424 12795
rect 16776 12764 16804 12795
rect 17420 12764 17448 12795
rect 17862 12792 17868 12804
rect 17920 12792 17926 12844
rect 14884 12736 17448 12764
rect 14884 12724 14890 12736
rect 9548 12668 10732 12696
rect 9548 12656 9554 12668
rect 11238 12656 11244 12708
rect 11296 12696 11302 12708
rect 11701 12699 11759 12705
rect 11701 12696 11713 12699
rect 11296 12668 11713 12696
rect 11296 12656 11302 12668
rect 11701 12665 11713 12668
rect 11747 12665 11759 12699
rect 11701 12659 11759 12665
rect 7392 12600 8156 12628
rect 8297 12631 8355 12637
rect 4755 12597 4767 12600
rect 4709 12591 4767 12597
rect 8297 12597 8309 12631
rect 8343 12628 8355 12631
rect 8570 12628 8576 12640
rect 8343 12600 8576 12628
rect 8343 12597 8355 12600
rect 8297 12591 8355 12597
rect 8570 12588 8576 12600
rect 8628 12588 8634 12640
rect 16666 12588 16672 12640
rect 16724 12628 16730 12640
rect 16761 12631 16819 12637
rect 16761 12628 16773 12631
rect 16724 12600 16773 12628
rect 16724 12588 16730 12600
rect 16761 12597 16773 12600
rect 16807 12597 16819 12631
rect 16761 12591 16819 12597
rect 16942 12588 16948 12640
rect 17000 12628 17006 12640
rect 17405 12631 17463 12637
rect 17405 12628 17417 12631
rect 17000 12600 17417 12628
rect 17000 12588 17006 12600
rect 17405 12597 17417 12600
rect 17451 12597 17463 12631
rect 17405 12591 17463 12597
rect 1104 12538 25852 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 12214 12538
rect 12266 12486 12278 12538
rect 12330 12486 12342 12538
rect 12394 12486 12406 12538
rect 12458 12486 12470 12538
rect 12522 12486 20214 12538
rect 20266 12486 20278 12538
rect 20330 12486 20342 12538
rect 20394 12486 20406 12538
rect 20458 12486 20470 12538
rect 20522 12486 25852 12538
rect 1104 12464 25852 12486
rect 10597 12427 10655 12433
rect 10597 12393 10609 12427
rect 10643 12424 10655 12427
rect 10870 12424 10876 12436
rect 10643 12396 10876 12424
rect 10643 12393 10655 12396
rect 10597 12387 10655 12393
rect 10870 12384 10876 12396
rect 10928 12384 10934 12436
rect 13449 12427 13507 12433
rect 13449 12424 13461 12427
rect 12406 12396 13461 12424
rect 7006 12356 7012 12368
rect 2700 12328 7012 12356
rect 2700 12232 2728 12328
rect 7006 12316 7012 12328
rect 7064 12316 7070 12368
rect 9766 12316 9772 12368
rect 9824 12356 9830 12368
rect 10134 12356 10140 12368
rect 9824 12328 10140 12356
rect 9824 12316 9830 12328
rect 10134 12316 10140 12328
rect 10192 12356 10198 12368
rect 12406 12356 12434 12396
rect 13449 12393 13461 12396
rect 13495 12393 13507 12427
rect 13449 12387 13507 12393
rect 16758 12384 16764 12436
rect 16816 12424 16822 12436
rect 17957 12427 18015 12433
rect 17957 12424 17969 12427
rect 16816 12396 17969 12424
rect 16816 12384 16822 12396
rect 17957 12393 17969 12396
rect 18003 12424 18015 12427
rect 18230 12424 18236 12436
rect 18003 12396 18236 12424
rect 18003 12393 18015 12396
rect 17957 12387 18015 12393
rect 18230 12384 18236 12396
rect 18288 12384 18294 12436
rect 10192 12328 12434 12356
rect 10192 12316 10198 12328
rect 4798 12248 4804 12300
rect 4856 12288 4862 12300
rect 4893 12291 4951 12297
rect 4893 12288 4905 12291
rect 4856 12260 4905 12288
rect 4856 12248 4862 12260
rect 4893 12257 4905 12260
rect 4939 12257 4951 12291
rect 7024 12288 7052 12316
rect 11790 12288 11796 12300
rect 7024 12260 11796 12288
rect 4893 12251 4951 12257
rect 11790 12248 11796 12260
rect 11848 12248 11854 12300
rect 15562 12248 15568 12300
rect 15620 12288 15626 12300
rect 16758 12288 16764 12300
rect 15620 12260 16764 12288
rect 15620 12248 15626 12260
rect 16758 12248 16764 12260
rect 16816 12248 16822 12300
rect 16850 12248 16856 12300
rect 16908 12288 16914 12300
rect 17494 12288 17500 12300
rect 16908 12260 17500 12288
rect 16908 12248 16914 12260
rect 17494 12248 17500 12260
rect 17552 12288 17558 12300
rect 19337 12291 19395 12297
rect 19337 12288 19349 12291
rect 17552 12260 19349 12288
rect 17552 12248 17558 12260
rect 19337 12257 19349 12260
rect 19383 12288 19395 12291
rect 19610 12288 19616 12300
rect 19383 12260 19616 12288
rect 19383 12257 19395 12260
rect 19337 12251 19395 12257
rect 19610 12248 19616 12260
rect 19668 12248 19674 12300
rect 2406 12180 2412 12232
rect 2464 12220 2470 12232
rect 2501 12223 2559 12229
rect 2501 12220 2513 12223
rect 2464 12192 2513 12220
rect 2464 12180 2470 12192
rect 2501 12189 2513 12192
rect 2547 12189 2559 12223
rect 2501 12183 2559 12189
rect 2682 12180 2688 12232
rect 2740 12180 2746 12232
rect 3418 12180 3424 12232
rect 3476 12220 3482 12232
rect 4187 12223 4245 12229
rect 4187 12220 4199 12223
rect 3476 12192 4199 12220
rect 3476 12180 3482 12192
rect 4187 12189 4199 12192
rect 4233 12189 4245 12223
rect 4187 12183 4245 12189
rect 4341 12223 4399 12229
rect 4341 12189 4353 12223
rect 4387 12189 4399 12223
rect 4341 12183 4399 12189
rect 4985 12223 5043 12229
rect 4985 12189 4997 12223
rect 5031 12189 5043 12223
rect 4985 12183 5043 12189
rect 5629 12223 5687 12229
rect 5629 12189 5641 12223
rect 5675 12220 5687 12223
rect 5994 12220 6000 12232
rect 5675 12192 6000 12220
rect 5675 12189 5687 12192
rect 5629 12183 5687 12189
rect 4356 12152 4384 12183
rect 4890 12152 4896 12164
rect 4356 12124 4896 12152
rect 4890 12112 4896 12124
rect 4948 12112 4954 12164
rect 5000 12152 5028 12183
rect 5994 12180 6000 12192
rect 6052 12180 6058 12232
rect 9674 12180 9680 12232
rect 9732 12180 9738 12232
rect 9861 12223 9919 12229
rect 9861 12189 9873 12223
rect 9907 12220 9919 12223
rect 9907 12192 10732 12220
rect 9907 12189 9919 12192
rect 9861 12183 9919 12189
rect 6270 12152 6276 12164
rect 5000 12124 6276 12152
rect 6270 12112 6276 12124
rect 6328 12112 6334 12164
rect 10704 12161 10732 12192
rect 11238 12180 11244 12232
rect 11296 12180 11302 12232
rect 11514 12180 11520 12232
rect 11572 12180 11578 12232
rect 13630 12180 13636 12232
rect 13688 12180 13694 12232
rect 14826 12180 14832 12232
rect 14884 12180 14890 12232
rect 15010 12180 15016 12232
rect 15068 12180 15074 12232
rect 17773 12223 17831 12229
rect 17773 12189 17785 12223
rect 17819 12189 17831 12223
rect 17773 12183 17831 12189
rect 10689 12155 10747 12161
rect 10689 12121 10701 12155
rect 10735 12121 10747 12155
rect 16942 12152 16948 12164
rect 16790 12124 16948 12152
rect 10689 12115 10747 12121
rect 2590 12044 2596 12096
rect 2648 12044 2654 12096
rect 3970 12044 3976 12096
rect 4028 12044 4034 12096
rect 5353 12087 5411 12093
rect 5353 12053 5365 12087
rect 5399 12084 5411 12087
rect 5534 12084 5540 12096
rect 5399 12056 5540 12084
rect 5399 12053 5411 12056
rect 5353 12047 5411 12053
rect 5534 12044 5540 12056
rect 5592 12044 5598 12096
rect 5810 12044 5816 12096
rect 5868 12044 5874 12096
rect 9766 12044 9772 12096
rect 9824 12044 9830 12096
rect 10704 12084 10732 12115
rect 16942 12112 16948 12124
rect 17000 12112 17006 12164
rect 17218 12112 17224 12164
rect 17276 12112 17282 12164
rect 11057 12087 11115 12093
rect 11057 12084 11069 12087
rect 10704 12056 11069 12084
rect 11057 12053 11069 12056
rect 11103 12053 11115 12087
rect 11057 12047 11115 12053
rect 11698 12044 11704 12096
rect 11756 12044 11762 12096
rect 14918 12044 14924 12096
rect 14976 12044 14982 12096
rect 15749 12087 15807 12093
rect 15749 12053 15761 12087
rect 15795 12084 15807 12087
rect 16574 12084 16580 12096
rect 15795 12056 16580 12084
rect 15795 12053 15807 12056
rect 15749 12047 15807 12053
rect 16574 12044 16580 12056
rect 16632 12044 16638 12096
rect 16850 12044 16856 12096
rect 16908 12084 16914 12096
rect 17788 12084 17816 12183
rect 18230 12180 18236 12232
rect 18288 12180 18294 12232
rect 18411 12223 18469 12229
rect 18411 12216 18423 12223
rect 18340 12189 18423 12216
rect 18457 12189 18469 12223
rect 18340 12188 18469 12189
rect 17862 12112 17868 12164
rect 17920 12152 17926 12164
rect 18340 12152 18368 12188
rect 18411 12183 18469 12188
rect 18506 12180 18512 12232
rect 18564 12220 18570 12232
rect 18693 12223 18751 12229
rect 18693 12220 18705 12223
rect 18564 12192 18705 12220
rect 18564 12180 18570 12192
rect 18693 12189 18705 12192
rect 18739 12189 18751 12223
rect 18693 12183 18751 12189
rect 18877 12223 18935 12229
rect 18877 12189 18889 12223
rect 18923 12189 18935 12223
rect 18877 12183 18935 12189
rect 18892 12152 18920 12183
rect 17920 12124 18920 12152
rect 17920 12112 17926 12124
rect 19518 12112 19524 12164
rect 19576 12152 19582 12164
rect 19613 12155 19671 12161
rect 19613 12152 19625 12155
rect 19576 12124 19625 12152
rect 19576 12112 19582 12124
rect 19613 12121 19625 12124
rect 19659 12121 19671 12155
rect 19613 12115 19671 12121
rect 19720 12124 20102 12152
rect 16908 12056 17816 12084
rect 16908 12044 16914 12056
rect 18322 12044 18328 12096
rect 18380 12044 18386 12096
rect 18785 12087 18843 12093
rect 18785 12053 18797 12087
rect 18831 12084 18843 12087
rect 19720 12084 19748 12124
rect 18831 12056 19748 12084
rect 18831 12053 18843 12056
rect 18785 12047 18843 12053
rect 20990 12044 20996 12096
rect 21048 12084 21054 12096
rect 21085 12087 21143 12093
rect 21085 12084 21097 12087
rect 21048 12056 21097 12084
rect 21048 12044 21054 12056
rect 21085 12053 21097 12056
rect 21131 12053 21143 12087
rect 21085 12047 21143 12053
rect 1104 11994 25852 12016
rect 1104 11942 8214 11994
rect 8266 11942 8278 11994
rect 8330 11942 8342 11994
rect 8394 11942 8406 11994
rect 8458 11942 8470 11994
rect 8522 11942 16214 11994
rect 16266 11942 16278 11994
rect 16330 11942 16342 11994
rect 16394 11942 16406 11994
rect 16458 11942 16470 11994
rect 16522 11942 24214 11994
rect 24266 11942 24278 11994
rect 24330 11942 24342 11994
rect 24394 11942 24406 11994
rect 24458 11942 24470 11994
rect 24522 11942 25852 11994
rect 1104 11920 25852 11942
rect 8570 11840 8576 11892
rect 8628 11840 8634 11892
rect 9861 11883 9919 11889
rect 9861 11849 9873 11883
rect 9907 11880 9919 11883
rect 10042 11880 10048 11892
rect 9907 11852 10048 11880
rect 9907 11849 9919 11852
rect 9861 11843 9919 11849
rect 10042 11840 10048 11852
rect 10100 11840 10106 11892
rect 10686 11840 10692 11892
rect 10744 11840 10750 11892
rect 11238 11840 11244 11892
rect 11296 11840 11302 11892
rect 11790 11840 11796 11892
rect 11848 11880 11854 11892
rect 13814 11880 13820 11892
rect 11848 11852 13820 11880
rect 11848 11840 11854 11852
rect 13814 11840 13820 11852
rect 13872 11840 13878 11892
rect 13998 11840 14004 11892
rect 14056 11840 14062 11892
rect 14274 11840 14280 11892
rect 14332 11880 14338 11892
rect 15933 11883 15991 11889
rect 15933 11880 15945 11883
rect 14332 11852 15945 11880
rect 14332 11840 14338 11852
rect 15933 11849 15945 11852
rect 15979 11849 15991 11883
rect 15933 11843 15991 11849
rect 17218 11840 17224 11892
rect 17276 11840 17282 11892
rect 20257 11883 20315 11889
rect 20257 11880 20269 11883
rect 18248 11852 20269 11880
rect 2590 11772 2596 11824
rect 2648 11772 2654 11824
rect 5718 11812 5724 11824
rect 5382 11784 5724 11812
rect 5718 11772 5724 11784
rect 5776 11772 5782 11824
rect 5810 11772 5816 11824
rect 5868 11772 5874 11824
rect 8389 11815 8447 11821
rect 8389 11781 8401 11815
rect 8435 11812 8447 11815
rect 8588 11812 8616 11840
rect 9766 11812 9772 11824
rect 8435 11784 8616 11812
rect 9614 11784 9772 11812
rect 8435 11781 8447 11784
rect 8389 11775 8447 11781
rect 9766 11772 9772 11784
rect 9824 11772 9830 11824
rect 11256 11812 11284 11840
rect 11701 11815 11759 11821
rect 11701 11812 11713 11815
rect 11256 11784 11713 11812
rect 11701 11781 11713 11784
rect 11747 11812 11759 11815
rect 12253 11815 12311 11821
rect 12253 11812 12265 11815
rect 11747 11784 12265 11812
rect 11747 11781 11759 11784
rect 11701 11775 11759 11781
rect 12253 11781 12265 11784
rect 12299 11781 12311 11815
rect 14016 11812 14044 11840
rect 14918 11812 14924 11824
rect 12253 11775 12311 11781
rect 13372 11784 14044 11812
rect 14858 11784 14924 11812
rect 3970 11744 3976 11756
rect 3931 11716 3976 11744
rect 3970 11704 3976 11716
rect 4028 11704 4034 11756
rect 4065 11747 4123 11753
rect 4065 11713 4077 11747
rect 4111 11744 4123 11747
rect 4522 11744 4528 11756
rect 4111 11716 4528 11744
rect 4111 11713 4123 11716
rect 4065 11707 4123 11713
rect 4522 11704 4528 11716
rect 4580 11704 4586 11756
rect 6089 11747 6147 11753
rect 6089 11713 6101 11747
rect 6135 11744 6147 11747
rect 6914 11744 6920 11756
rect 6135 11716 6920 11744
rect 6135 11713 6147 11716
rect 6089 11707 6147 11713
rect 6914 11704 6920 11716
rect 6972 11744 6978 11756
rect 7834 11744 7840 11756
rect 6972 11716 7840 11744
rect 6972 11704 6978 11716
rect 7834 11704 7840 11716
rect 7892 11744 7898 11756
rect 8113 11747 8171 11753
rect 8113 11744 8125 11747
rect 7892 11716 8125 11744
rect 7892 11704 7898 11716
rect 8113 11713 8125 11716
rect 8159 11713 8171 11747
rect 8113 11707 8171 11713
rect 10318 11704 10324 11756
rect 10376 11744 10382 11756
rect 13372 11753 13400 11784
rect 14918 11772 14924 11784
rect 14976 11772 14982 11824
rect 18248 11812 18276 11852
rect 20257 11849 20269 11852
rect 20303 11849 20315 11883
rect 20257 11843 20315 11849
rect 15028 11784 18276 11812
rect 10413 11747 10471 11753
rect 10413 11744 10425 11747
rect 10376 11716 10425 11744
rect 10376 11704 10382 11716
rect 10413 11713 10425 11716
rect 10459 11713 10471 11747
rect 11057 11747 11115 11753
rect 11057 11744 11069 11747
rect 10413 11707 10471 11713
rect 10520 11716 11069 11744
rect 1486 11636 1492 11688
rect 1544 11676 1550 11688
rect 1673 11679 1731 11685
rect 1673 11676 1685 11679
rect 1544 11648 1685 11676
rect 1544 11636 1550 11648
rect 1673 11645 1685 11648
rect 1719 11645 1731 11679
rect 1673 11639 1731 11645
rect 1946 11636 1952 11688
rect 2004 11636 2010 11688
rect 2406 11636 2412 11688
rect 2464 11676 2470 11688
rect 6822 11676 6828 11688
rect 2464 11648 6828 11676
rect 2464 11636 2470 11648
rect 6822 11636 6828 11648
rect 6880 11636 6886 11688
rect 10520 11676 10548 11716
rect 11057 11713 11069 11716
rect 11103 11713 11115 11747
rect 11057 11707 11115 11713
rect 11241 11747 11299 11753
rect 11241 11713 11253 11747
rect 11287 11713 11299 11747
rect 11241 11707 11299 11713
rect 13357 11747 13415 11753
rect 13357 11713 13369 11747
rect 13403 11713 13415 11747
rect 13357 11707 13415 11713
rect 6932 11648 10548 11676
rect 10781 11679 10839 11685
rect 3697 11611 3755 11617
rect 3697 11577 3709 11611
rect 3743 11608 3755 11611
rect 4614 11608 4620 11620
rect 3743 11580 4620 11608
rect 3743 11577 3755 11580
rect 3697 11571 3755 11577
rect 4614 11568 4620 11580
rect 4672 11568 4678 11620
rect 6730 11568 6736 11620
rect 6788 11608 6794 11620
rect 6932 11608 6960 11648
rect 10781 11645 10793 11679
rect 10827 11676 10839 11679
rect 11256 11676 11284 11707
rect 13633 11679 13691 11685
rect 13633 11676 13645 11679
rect 10827 11648 11284 11676
rect 13464 11648 13645 11676
rect 10827 11645 10839 11648
rect 10781 11639 10839 11645
rect 6788 11580 6960 11608
rect 6788 11568 6794 11580
rect 11422 11568 11428 11620
rect 11480 11608 11486 11620
rect 12437 11611 12495 11617
rect 11480 11580 11928 11608
rect 11480 11568 11486 11580
rect 3418 11500 3424 11552
rect 3476 11500 3482 11552
rect 4062 11500 4068 11552
rect 4120 11540 4126 11552
rect 4341 11543 4399 11549
rect 4341 11540 4353 11543
rect 4120 11512 4353 11540
rect 4120 11500 4126 11512
rect 4341 11509 4353 11512
rect 4387 11509 4399 11543
rect 4341 11503 4399 11509
rect 9950 11500 9956 11552
rect 10008 11540 10014 11552
rect 10229 11543 10287 11549
rect 10229 11540 10241 11543
rect 10008 11512 10241 11540
rect 10008 11500 10014 11512
rect 10229 11509 10241 11512
rect 10275 11509 10287 11543
rect 11900 11540 11928 11580
rect 12437 11577 12449 11611
rect 12483 11608 12495 11611
rect 12802 11608 12808 11620
rect 12483 11580 12808 11608
rect 12483 11577 12495 11580
rect 12437 11571 12495 11577
rect 12802 11568 12808 11580
rect 12860 11568 12866 11620
rect 13354 11568 13360 11620
rect 13412 11608 13418 11620
rect 13464 11608 13492 11648
rect 13633 11645 13645 11648
rect 13679 11645 13691 11679
rect 13633 11639 13691 11645
rect 13412 11580 13492 11608
rect 13412 11568 13418 11580
rect 15028 11540 15056 11784
rect 18322 11772 18328 11824
rect 18380 11812 18386 11824
rect 18380 11784 18538 11812
rect 18380 11772 18386 11784
rect 16025 11747 16083 11753
rect 16025 11713 16037 11747
rect 16071 11744 16083 11747
rect 16574 11744 16580 11756
rect 16071 11716 16580 11744
rect 16071 11713 16083 11716
rect 16025 11707 16083 11713
rect 16574 11704 16580 11716
rect 16632 11704 16638 11756
rect 16758 11704 16764 11756
rect 16816 11704 16822 11756
rect 17405 11747 17463 11753
rect 17405 11713 17417 11747
rect 17451 11713 17463 11747
rect 17405 11707 17463 11713
rect 15841 11679 15899 11685
rect 15841 11645 15853 11679
rect 15887 11645 15899 11679
rect 17420 11676 17448 11707
rect 17494 11704 17500 11756
rect 17552 11744 17558 11756
rect 17773 11747 17831 11753
rect 17773 11744 17785 11747
rect 17552 11716 17785 11744
rect 17552 11704 17558 11716
rect 17773 11713 17785 11716
rect 17819 11713 17831 11747
rect 17773 11707 17831 11713
rect 20165 11747 20223 11753
rect 20165 11713 20177 11747
rect 20211 11744 20223 11747
rect 20990 11744 20996 11756
rect 20211 11716 20996 11744
rect 20211 11713 20223 11716
rect 20165 11707 20223 11713
rect 20990 11704 20996 11716
rect 21048 11704 21054 11756
rect 15841 11639 15899 11645
rect 16546 11648 17448 11676
rect 15856 11608 15884 11639
rect 16022 11608 16028 11620
rect 15856 11580 16028 11608
rect 16022 11568 16028 11580
rect 16080 11568 16086 11620
rect 16393 11611 16451 11617
rect 16393 11577 16405 11611
rect 16439 11608 16451 11611
rect 16546 11608 16574 11648
rect 18046 11636 18052 11688
rect 18104 11636 18110 11688
rect 19978 11636 19984 11688
rect 20036 11676 20042 11688
rect 20349 11679 20407 11685
rect 20349 11676 20361 11679
rect 20036 11648 20361 11676
rect 20036 11636 20042 11648
rect 20349 11645 20361 11648
rect 20395 11645 20407 11679
rect 20349 11639 20407 11645
rect 16439 11580 16574 11608
rect 16439 11577 16451 11580
rect 16393 11571 16451 11577
rect 19058 11568 19064 11620
rect 19116 11608 19122 11620
rect 19521 11611 19579 11617
rect 19521 11608 19533 11611
rect 19116 11580 19533 11608
rect 19116 11568 19122 11580
rect 19521 11577 19533 11580
rect 19567 11608 19579 11611
rect 22646 11608 22652 11620
rect 19567 11580 22652 11608
rect 19567 11577 19579 11580
rect 19521 11571 19579 11577
rect 22646 11568 22652 11580
rect 22704 11568 22710 11620
rect 11900 11512 15056 11540
rect 10229 11503 10287 11509
rect 15102 11500 15108 11552
rect 15160 11500 15166 11552
rect 16942 11500 16948 11552
rect 17000 11500 17006 11552
rect 19794 11500 19800 11552
rect 19852 11500 19858 11552
rect 1104 11450 25852 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 12214 11450
rect 12266 11398 12278 11450
rect 12330 11398 12342 11450
rect 12394 11398 12406 11450
rect 12458 11398 12470 11450
rect 12522 11398 20214 11450
rect 20266 11398 20278 11450
rect 20330 11398 20342 11450
rect 20394 11398 20406 11450
rect 20458 11398 20470 11450
rect 20522 11398 25852 11450
rect 1104 11376 25852 11398
rect 1946 11296 1952 11348
rect 2004 11336 2010 11348
rect 2225 11339 2283 11345
rect 2225 11336 2237 11339
rect 2004 11308 2237 11336
rect 2004 11296 2010 11308
rect 2225 11305 2237 11308
rect 2271 11305 2283 11339
rect 2225 11299 2283 11305
rect 3344 11308 4752 11336
rect 2777 11271 2835 11277
rect 2777 11237 2789 11271
rect 2823 11237 2835 11271
rect 2777 11231 2835 11237
rect 2409 11135 2467 11141
rect 2409 11101 2421 11135
rect 2455 11132 2467 11135
rect 2792 11132 2820 11231
rect 3344 11212 3372 11308
rect 3970 11228 3976 11280
rect 4028 11268 4034 11280
rect 4028 11240 4660 11268
rect 4028 11228 4034 11240
rect 3326 11160 3332 11212
rect 3384 11160 3390 11212
rect 4433 11203 4491 11209
rect 4433 11169 4445 11203
rect 4479 11169 4491 11203
rect 4433 11163 4491 11169
rect 2455 11104 2820 11132
rect 3145 11135 3203 11141
rect 2455 11101 2467 11104
rect 2409 11095 2467 11101
rect 3145 11101 3157 11135
rect 3191 11132 3203 11135
rect 3418 11132 3424 11144
rect 3191 11104 3424 11132
rect 3191 11101 3203 11104
rect 3145 11095 3203 11101
rect 3418 11092 3424 11104
rect 3476 11132 3482 11144
rect 3970 11132 3976 11144
rect 3476 11104 3976 11132
rect 3476 11092 3482 11104
rect 3970 11092 3976 11104
rect 4028 11132 4034 11144
rect 4448 11132 4476 11163
rect 4028 11104 4476 11132
rect 4525 11135 4583 11141
rect 4028 11092 4034 11104
rect 4525 11101 4537 11135
rect 4571 11101 4583 11135
rect 4632 11132 4660 11240
rect 4724 11200 4752 11308
rect 4798 11296 4804 11348
rect 4856 11296 4862 11348
rect 5994 11296 6000 11348
rect 6052 11296 6058 11348
rect 6270 11296 6276 11348
rect 6328 11296 6334 11348
rect 9950 11345 9956 11348
rect 9940 11339 9956 11345
rect 9940 11305 9952 11339
rect 9940 11299 9956 11305
rect 9950 11296 9956 11299
rect 10008 11296 10014 11348
rect 11422 11296 11428 11348
rect 11480 11296 11486 11348
rect 11698 11296 11704 11348
rect 11756 11336 11762 11348
rect 11958 11339 12016 11345
rect 11958 11336 11970 11339
rect 11756 11308 11970 11336
rect 11756 11296 11762 11308
rect 11958 11305 11970 11308
rect 12004 11305 12016 11339
rect 11958 11299 12016 11305
rect 12158 11296 12164 11348
rect 12216 11336 12222 11348
rect 14274 11336 14280 11348
rect 12216 11308 14280 11336
rect 12216 11296 12222 11308
rect 14274 11296 14280 11308
rect 14332 11296 14338 11348
rect 14826 11296 14832 11348
rect 14884 11296 14890 11348
rect 17957 11339 18015 11345
rect 17957 11305 17969 11339
rect 18003 11336 18015 11339
rect 18046 11336 18052 11348
rect 18003 11308 18052 11336
rect 18003 11305 18015 11308
rect 17957 11299 18015 11305
rect 18046 11296 18052 11308
rect 18104 11296 18110 11348
rect 19518 11296 19524 11348
rect 19576 11296 19582 11348
rect 21913 11339 21971 11345
rect 21913 11305 21925 11339
rect 21959 11336 21971 11339
rect 22278 11336 22284 11348
rect 21959 11308 22284 11336
rect 21959 11305 21971 11308
rect 21913 11299 21971 11305
rect 22278 11296 22284 11308
rect 22336 11296 22342 11348
rect 5368 11240 5672 11268
rect 5368 11209 5396 11240
rect 5353 11203 5411 11209
rect 5353 11200 5365 11203
rect 4724 11172 5365 11200
rect 5353 11169 5365 11172
rect 5399 11169 5411 11203
rect 5353 11163 5411 11169
rect 5534 11160 5540 11212
rect 5592 11160 5598 11212
rect 5644 11200 5672 11240
rect 5718 11228 5724 11280
rect 5776 11268 5782 11280
rect 7009 11271 7067 11277
rect 7009 11268 7021 11271
rect 5776 11240 7021 11268
rect 5776 11228 5782 11240
rect 7009 11237 7021 11240
rect 7055 11237 7067 11271
rect 7009 11231 7067 11237
rect 7653 11271 7711 11277
rect 7653 11237 7665 11271
rect 7699 11268 7711 11271
rect 7742 11268 7748 11280
rect 7699 11240 7748 11268
rect 7699 11237 7711 11240
rect 7653 11231 7711 11237
rect 7742 11228 7748 11240
rect 7800 11228 7806 11280
rect 7834 11228 7840 11280
rect 7892 11228 7898 11280
rect 14369 11271 14427 11277
rect 14369 11237 14381 11271
rect 14415 11268 14427 11271
rect 15562 11268 15568 11280
rect 14415 11240 15568 11268
rect 14415 11237 14427 11240
rect 14369 11231 14427 11237
rect 15562 11228 15568 11240
rect 15620 11228 15626 11280
rect 18233 11271 18291 11277
rect 18233 11237 18245 11271
rect 18279 11237 18291 11271
rect 18233 11231 18291 11237
rect 20533 11271 20591 11277
rect 20533 11237 20545 11271
rect 20579 11237 20591 11271
rect 20533 11231 20591 11237
rect 22189 11271 22247 11277
rect 22189 11237 22201 11271
rect 22235 11237 22247 11271
rect 22189 11231 22247 11237
rect 7374 11200 7380 11212
rect 5644 11172 7380 11200
rect 7374 11160 7380 11172
rect 7432 11160 7438 11212
rect 7852 11200 7880 11228
rect 9677 11203 9735 11209
rect 9677 11200 9689 11203
rect 7852 11172 9689 11200
rect 9677 11169 9689 11172
rect 9723 11200 9735 11203
rect 10410 11200 10416 11212
rect 9723 11172 10416 11200
rect 9723 11169 9735 11172
rect 9677 11163 9735 11169
rect 10410 11160 10416 11172
rect 10468 11200 10474 11212
rect 11701 11203 11759 11209
rect 11701 11200 11713 11203
rect 10468 11172 11713 11200
rect 10468 11160 10474 11172
rect 11701 11169 11713 11172
rect 11747 11200 11759 11203
rect 13998 11200 14004 11212
rect 11747 11172 14004 11200
rect 11747 11169 11759 11172
rect 11701 11163 11759 11169
rect 13998 11160 14004 11172
rect 14056 11160 14062 11212
rect 16942 11160 16948 11212
rect 17000 11160 17006 11212
rect 17221 11203 17279 11209
rect 17221 11169 17233 11203
rect 17267 11200 17279 11203
rect 17494 11200 17500 11212
rect 17267 11172 17500 11200
rect 17267 11169 17279 11172
rect 17221 11163 17279 11169
rect 17494 11160 17500 11172
rect 17552 11160 17558 11212
rect 6457 11135 6515 11141
rect 6457 11132 6469 11135
rect 4632 11104 6469 11132
rect 4525 11095 4583 11101
rect 6457 11101 6469 11104
rect 6503 11101 6515 11135
rect 6457 11095 6515 11101
rect 4062 11024 4068 11076
rect 4120 11064 4126 11076
rect 4540 11064 4568 11095
rect 6546 11092 6552 11144
rect 6604 11092 6610 11144
rect 6822 11092 6828 11144
rect 6880 11092 6886 11144
rect 7006 11092 7012 11144
rect 7064 11092 7070 11144
rect 7837 11135 7895 11141
rect 7837 11101 7849 11135
rect 7883 11132 7895 11135
rect 7926 11132 7932 11144
rect 7883 11104 7932 11132
rect 7883 11101 7895 11104
rect 7837 11095 7895 11101
rect 7926 11092 7932 11104
rect 7984 11092 7990 11144
rect 8297 11135 8355 11141
rect 8297 11101 8309 11135
rect 8343 11132 8355 11135
rect 9030 11132 9036 11144
rect 8343 11104 9036 11132
rect 8343 11101 8355 11104
rect 8297 11095 8355 11101
rect 9030 11092 9036 11104
rect 9088 11092 9094 11144
rect 9217 11135 9275 11141
rect 9217 11101 9229 11135
rect 9263 11101 9275 11135
rect 9217 11095 9275 11101
rect 9401 11135 9459 11141
rect 9401 11101 9413 11135
rect 9447 11101 9459 11135
rect 9401 11095 9459 11101
rect 4120 11036 4568 11064
rect 4120 11024 4126 11036
rect 3234 10956 3240 11008
rect 3292 10956 3298 11008
rect 4540 10996 4568 11036
rect 4706 11024 4712 11076
rect 4764 11064 4770 11076
rect 6273 11067 6331 11073
rect 6273 11064 6285 11067
rect 4764 11036 6285 11064
rect 4764 11024 4770 11036
rect 6273 11033 6285 11036
rect 6319 11033 6331 11067
rect 6273 11027 6331 11033
rect 4798 10996 4804 11008
rect 4540 10968 4804 10996
rect 4798 10956 4804 10968
rect 4856 10996 4862 11008
rect 5629 10999 5687 11005
rect 5629 10996 5641 10999
rect 4856 10968 5641 10996
rect 4856 10956 4862 10968
rect 5629 10965 5641 10968
rect 5675 10965 5687 10999
rect 5629 10959 5687 10965
rect 8110 10956 8116 11008
rect 8168 10956 8174 11008
rect 9232 10996 9260 11095
rect 9306 11024 9312 11076
rect 9364 11024 9370 11076
rect 9416 11064 9444 11095
rect 11054 11092 11060 11144
rect 11112 11092 11118 11144
rect 13630 11092 13636 11144
rect 13688 11132 13694 11144
rect 14185 11135 14243 11141
rect 14185 11132 14197 11135
rect 13688 11104 14197 11132
rect 13688 11092 13694 11104
rect 14185 11101 14197 11104
rect 14231 11101 14243 11135
rect 14185 11095 14243 11101
rect 17773 11135 17831 11141
rect 17773 11101 17785 11135
rect 17819 11132 17831 11135
rect 18248 11132 18276 11231
rect 18877 11203 18935 11209
rect 18877 11169 18889 11203
rect 18923 11200 18935 11203
rect 19978 11200 19984 11212
rect 18923 11172 19984 11200
rect 18923 11169 18935 11172
rect 18877 11163 18935 11169
rect 19978 11160 19984 11172
rect 20036 11160 20042 11212
rect 17819 11104 18276 11132
rect 18601 11135 18659 11141
rect 17819 11101 17831 11104
rect 17773 11095 17831 11101
rect 18601 11101 18613 11135
rect 18647 11132 18659 11135
rect 19058 11132 19064 11144
rect 18647 11104 19064 11132
rect 18647 11101 18659 11104
rect 18601 11095 18659 11101
rect 19058 11092 19064 11104
rect 19116 11092 19122 11144
rect 19337 11135 19395 11141
rect 19337 11101 19349 11135
rect 19383 11132 19395 11135
rect 19794 11132 19800 11144
rect 19383 11104 19800 11132
rect 19383 11101 19395 11104
rect 19337 11095 19395 11101
rect 19794 11092 19800 11104
rect 19852 11092 19858 11144
rect 20073 11135 20131 11141
rect 20073 11101 20085 11135
rect 20119 11132 20131 11135
rect 20548 11132 20576 11231
rect 20990 11160 20996 11212
rect 21048 11160 21054 11212
rect 21177 11203 21235 11209
rect 21177 11169 21189 11203
rect 21223 11200 21235 11203
rect 21223 11172 21312 11200
rect 21223 11169 21235 11172
rect 21177 11163 21235 11169
rect 20119 11104 20576 11132
rect 20119 11101 20131 11104
rect 20073 11095 20131 11101
rect 9416 11036 9996 11064
rect 9858 10996 9864 11008
rect 9232 10968 9864 10996
rect 9858 10956 9864 10968
rect 9916 10956 9922 11008
rect 9968 10996 9996 11036
rect 12618 11024 12624 11076
rect 12676 11024 12682 11076
rect 13814 11024 13820 11076
rect 13872 11064 13878 11076
rect 14734 11064 14740 11076
rect 13872 11036 14740 11064
rect 13872 11024 13878 11036
rect 14734 11024 14740 11036
rect 14792 11024 14798 11076
rect 16666 11064 16672 11076
rect 16514 11036 16672 11064
rect 16666 11024 16672 11036
rect 16724 11024 16730 11076
rect 18046 11024 18052 11076
rect 18104 11064 18110 11076
rect 18693 11067 18751 11073
rect 18693 11064 18705 11067
rect 18104 11036 18705 11064
rect 18104 11024 18110 11036
rect 18693 11033 18705 11036
rect 18739 11033 18751 11067
rect 21284 11064 21312 11172
rect 21729 11135 21787 11141
rect 21729 11101 21741 11135
rect 21775 11132 21787 11135
rect 22204 11132 22232 11231
rect 22646 11160 22652 11212
rect 22704 11160 22710 11212
rect 22833 11203 22891 11209
rect 22833 11169 22845 11203
rect 22879 11200 22891 11203
rect 23382 11200 23388 11212
rect 22879 11172 23388 11200
rect 22879 11169 22891 11172
rect 22833 11163 22891 11169
rect 22848 11132 22876 11163
rect 23382 11160 23388 11172
rect 23440 11160 23446 11212
rect 21775 11104 22232 11132
rect 22296 11104 22876 11132
rect 21775 11101 21787 11104
rect 21729 11095 21787 11101
rect 22296 11064 22324 11104
rect 18693 11027 18751 11033
rect 19996 11036 22324 11064
rect 22557 11067 22615 11073
rect 10042 10996 10048 11008
rect 9968 10968 10048 10996
rect 10042 10956 10048 10968
rect 10100 10996 10106 11008
rect 11238 10996 11244 11008
rect 10100 10968 11244 10996
rect 10100 10956 10106 10968
rect 11238 10956 11244 10968
rect 11296 10956 11302 11008
rect 12710 10956 12716 11008
rect 12768 10996 12774 11008
rect 13449 10999 13507 11005
rect 13449 10996 13461 10999
rect 12768 10968 13461 10996
rect 12768 10956 12774 10968
rect 13449 10965 13461 10968
rect 13495 10996 13507 10999
rect 13722 10996 13728 11008
rect 13495 10968 13728 10996
rect 13495 10965 13507 10968
rect 13449 10959 13507 10965
rect 13722 10956 13728 10968
rect 13780 10956 13786 11008
rect 15470 10956 15476 11008
rect 15528 10956 15534 11008
rect 18230 10956 18236 11008
rect 18288 10996 18294 11008
rect 19996 10996 20024 11036
rect 22557 11033 22569 11067
rect 22603 11064 22615 11067
rect 23842 11064 23848 11076
rect 22603 11036 23848 11064
rect 22603 11033 22615 11036
rect 22557 11027 22615 11033
rect 23842 11024 23848 11036
rect 23900 11024 23906 11076
rect 18288 10968 20024 10996
rect 18288 10956 18294 10968
rect 20070 10956 20076 11008
rect 20128 10996 20134 11008
rect 20257 10999 20315 11005
rect 20257 10996 20269 10999
rect 20128 10968 20269 10996
rect 20128 10956 20134 10968
rect 20257 10965 20269 10968
rect 20303 10965 20315 10999
rect 20257 10959 20315 10965
rect 20901 10999 20959 11005
rect 20901 10965 20913 10999
rect 20947 10996 20959 10999
rect 21910 10996 21916 11008
rect 20947 10968 21916 10996
rect 20947 10965 20959 10968
rect 20901 10959 20959 10965
rect 21910 10956 21916 10968
rect 21968 10956 21974 11008
rect 1104 10906 25852 10928
rect 1104 10854 8214 10906
rect 8266 10854 8278 10906
rect 8330 10854 8342 10906
rect 8394 10854 8406 10906
rect 8458 10854 8470 10906
rect 8522 10854 16214 10906
rect 16266 10854 16278 10906
rect 16330 10854 16342 10906
rect 16394 10854 16406 10906
rect 16458 10854 16470 10906
rect 16522 10854 24214 10906
rect 24266 10854 24278 10906
rect 24330 10854 24342 10906
rect 24394 10854 24406 10906
rect 24458 10854 24470 10906
rect 24522 10854 25852 10906
rect 1104 10832 25852 10854
rect 3234 10752 3240 10804
rect 3292 10792 3298 10804
rect 3881 10795 3939 10801
rect 3881 10792 3893 10795
rect 3292 10764 3893 10792
rect 3292 10752 3298 10764
rect 3881 10761 3893 10764
rect 3927 10761 3939 10795
rect 3881 10755 3939 10761
rect 4706 10752 4712 10804
rect 4764 10752 4770 10804
rect 4982 10752 4988 10804
rect 5040 10792 5046 10804
rect 6914 10792 6920 10804
rect 5040 10764 6920 10792
rect 5040 10752 5046 10764
rect 6914 10752 6920 10764
rect 6972 10752 6978 10804
rect 7374 10752 7380 10804
rect 7432 10752 7438 10804
rect 8018 10792 8024 10804
rect 7576 10764 8024 10792
rect 1302 10684 1308 10736
rect 1360 10724 1366 10736
rect 3605 10727 3663 10733
rect 1360 10696 3280 10724
rect 1360 10684 1366 10696
rect 2406 10616 2412 10668
rect 2464 10616 2470 10668
rect 2593 10659 2651 10665
rect 2593 10625 2605 10659
rect 2639 10656 2651 10659
rect 2682 10656 2688 10668
rect 2639 10628 2688 10656
rect 2639 10625 2651 10628
rect 2593 10619 2651 10625
rect 2682 10616 2688 10628
rect 2740 10616 2746 10668
rect 3252 10665 3280 10696
rect 3605 10693 3617 10727
rect 3651 10724 3663 10727
rect 6638 10724 6644 10736
rect 3651 10696 6644 10724
rect 3651 10693 3663 10696
rect 3605 10687 3663 10693
rect 6638 10684 6644 10696
rect 6696 10684 6702 10736
rect 3237 10659 3295 10665
rect 3237 10625 3249 10659
rect 3283 10625 3295 10659
rect 3237 10619 3295 10625
rect 3391 10659 3449 10665
rect 3391 10625 3403 10659
rect 3437 10656 3449 10659
rect 3970 10656 3976 10668
rect 3437 10628 3976 10656
rect 3437 10625 3449 10628
rect 3391 10619 3449 10625
rect 3252 10588 3280 10619
rect 3970 10616 3976 10628
rect 4028 10616 4034 10668
rect 4249 10659 4307 10665
rect 4249 10625 4261 10659
rect 4295 10656 4307 10659
rect 4614 10656 4620 10668
rect 4295 10628 4620 10656
rect 4295 10625 4307 10628
rect 4249 10619 4307 10625
rect 4614 10616 4620 10628
rect 4672 10616 4678 10668
rect 5720 10659 5778 10665
rect 5720 10625 5732 10659
rect 5766 10625 5778 10659
rect 5720 10619 5778 10625
rect 4062 10588 4068 10600
rect 3252 10560 4068 10588
rect 4062 10548 4068 10560
rect 4120 10548 4126 10600
rect 4341 10591 4399 10597
rect 4341 10557 4353 10591
rect 4387 10588 4399 10591
rect 5169 10591 5227 10597
rect 4387 10560 5120 10588
rect 4387 10557 4399 10560
rect 4341 10551 4399 10557
rect 3234 10480 3240 10532
rect 3292 10520 3298 10532
rect 4801 10523 4859 10529
rect 4801 10520 4813 10523
rect 3292 10492 4813 10520
rect 3292 10480 3298 10492
rect 4801 10489 4813 10492
rect 4847 10489 4859 10523
rect 5092 10520 5120 10560
rect 5169 10557 5181 10591
rect 5215 10588 5227 10591
rect 5534 10588 5540 10600
rect 5215 10560 5540 10588
rect 5215 10557 5227 10560
rect 5169 10551 5227 10557
rect 5534 10548 5540 10560
rect 5592 10548 5598 10600
rect 5736 10588 5764 10619
rect 5810 10616 5816 10668
rect 5868 10616 5874 10668
rect 6086 10616 6092 10668
rect 6144 10656 6150 10668
rect 7576 10665 7604 10764
rect 8018 10752 8024 10764
rect 8076 10792 8082 10804
rect 8076 10764 10088 10792
rect 8076 10752 8082 10764
rect 8110 10684 8116 10736
rect 8168 10684 8174 10736
rect 9953 10727 10011 10733
rect 9953 10724 9965 10727
rect 9338 10696 9965 10724
rect 9953 10693 9965 10696
rect 9999 10693 10011 10727
rect 10060 10724 10088 10764
rect 10318 10752 10324 10804
rect 10376 10792 10382 10804
rect 10413 10795 10471 10801
rect 10413 10792 10425 10795
rect 10376 10764 10425 10792
rect 10376 10752 10382 10764
rect 10413 10761 10425 10764
rect 10459 10761 10471 10795
rect 10413 10755 10471 10761
rect 10873 10795 10931 10801
rect 10873 10761 10885 10795
rect 10919 10792 10931 10795
rect 11422 10792 11428 10804
rect 10919 10764 11428 10792
rect 10919 10761 10931 10764
rect 10873 10755 10931 10761
rect 11422 10752 11428 10764
rect 11480 10752 11486 10804
rect 11514 10752 11520 10804
rect 11572 10792 11578 10804
rect 11609 10795 11667 10801
rect 11609 10792 11621 10795
rect 11572 10764 11621 10792
rect 11572 10752 11578 10764
rect 11609 10761 11621 10764
rect 11655 10761 11667 10795
rect 11609 10755 11667 10761
rect 12069 10795 12127 10801
rect 12069 10761 12081 10795
rect 12115 10792 12127 10795
rect 12710 10792 12716 10804
rect 12115 10764 12716 10792
rect 12115 10761 12127 10764
rect 12069 10755 12127 10761
rect 12710 10752 12716 10764
rect 12768 10752 12774 10804
rect 13354 10752 13360 10804
rect 13412 10752 13418 10804
rect 13633 10795 13691 10801
rect 13633 10761 13645 10795
rect 13679 10761 13691 10795
rect 13633 10755 13691 10761
rect 12342 10724 12348 10736
rect 10060 10696 12348 10724
rect 9953 10687 10011 10693
rect 12342 10684 12348 10696
rect 12400 10684 12406 10736
rect 12621 10727 12679 10733
rect 12621 10693 12633 10727
rect 12667 10724 12679 10727
rect 12894 10724 12900 10736
rect 12667 10696 12900 10724
rect 12667 10693 12679 10696
rect 12621 10687 12679 10693
rect 12894 10684 12900 10696
rect 12952 10684 12958 10736
rect 6733 10659 6791 10665
rect 6733 10656 6745 10659
rect 6144 10628 6745 10656
rect 6144 10616 6150 10628
rect 6733 10625 6745 10628
rect 6779 10625 6791 10659
rect 6733 10619 6791 10625
rect 7561 10659 7619 10665
rect 7561 10625 7573 10659
rect 7607 10625 7619 10659
rect 7561 10619 7619 10625
rect 7834 10616 7840 10668
rect 7892 10616 7898 10668
rect 9858 10616 9864 10668
rect 9916 10616 9922 10668
rect 10042 10616 10048 10668
rect 10100 10616 10106 10668
rect 10778 10616 10784 10668
rect 10836 10616 10842 10668
rect 11330 10616 11336 10668
rect 11388 10656 11394 10668
rect 11977 10659 12035 10665
rect 11977 10656 11989 10659
rect 11388 10628 11989 10656
rect 11388 10616 11394 10628
rect 11977 10625 11989 10628
rect 12023 10625 12035 10659
rect 11977 10619 12035 10625
rect 12084 10628 12296 10656
rect 6178 10588 6184 10600
rect 5736 10560 6184 10588
rect 6178 10548 6184 10560
rect 6236 10548 6242 10600
rect 6454 10548 6460 10600
rect 6512 10548 6518 10600
rect 10318 10548 10324 10600
rect 10376 10588 10382 10600
rect 11057 10591 11115 10597
rect 11057 10588 11069 10591
rect 10376 10560 11069 10588
rect 10376 10548 10382 10560
rect 11057 10557 11069 10560
rect 11103 10588 11115 10591
rect 12084 10588 12112 10628
rect 12268 10597 12296 10628
rect 12710 10616 12716 10668
rect 12768 10656 12774 10668
rect 12805 10659 12863 10665
rect 12805 10656 12817 10659
rect 12768 10628 12817 10656
rect 12768 10616 12774 10628
rect 12805 10625 12817 10628
rect 12851 10625 12863 10659
rect 12805 10619 12863 10625
rect 13173 10659 13231 10665
rect 13173 10625 13185 10659
rect 13219 10656 13231 10659
rect 13648 10656 13676 10755
rect 13722 10752 13728 10804
rect 13780 10792 13786 10804
rect 15565 10795 15623 10801
rect 15565 10792 15577 10795
rect 13780 10764 15577 10792
rect 13780 10752 13786 10764
rect 15565 10761 15577 10764
rect 15611 10761 15623 10795
rect 15565 10755 15623 10761
rect 16025 10795 16083 10801
rect 16025 10761 16037 10795
rect 16071 10792 16083 10795
rect 16758 10792 16764 10804
rect 16071 10764 16764 10792
rect 16071 10761 16083 10764
rect 16025 10755 16083 10761
rect 16758 10752 16764 10764
rect 16816 10752 16822 10804
rect 22554 10792 22560 10804
rect 21008 10764 22560 10792
rect 14001 10727 14059 10733
rect 14001 10693 14013 10727
rect 14047 10724 14059 10727
rect 15102 10724 15108 10736
rect 14047 10696 15108 10724
rect 14047 10693 14059 10696
rect 14001 10687 14059 10693
rect 15102 10684 15108 10696
rect 15160 10684 15166 10736
rect 15286 10684 15292 10736
rect 15344 10724 15350 10736
rect 18046 10724 18052 10736
rect 15344 10696 18052 10724
rect 15344 10684 15350 10696
rect 18046 10684 18052 10696
rect 18104 10684 18110 10736
rect 13219 10628 13676 10656
rect 14829 10659 14887 10665
rect 13219 10625 13231 10628
rect 13173 10619 13231 10625
rect 14829 10625 14841 10659
rect 14875 10656 14887 10659
rect 14918 10656 14924 10668
rect 14875 10628 14924 10656
rect 14875 10625 14887 10628
rect 14829 10619 14887 10625
rect 14918 10616 14924 10628
rect 14976 10616 14982 10668
rect 15470 10616 15476 10668
rect 15528 10656 15534 10668
rect 15657 10659 15715 10665
rect 15657 10656 15669 10659
rect 15528 10628 15669 10656
rect 15528 10616 15534 10628
rect 15657 10625 15669 10628
rect 15703 10656 15715 10659
rect 16114 10656 16120 10668
rect 15703 10628 16120 10656
rect 15703 10625 15715 10628
rect 15657 10619 15715 10625
rect 16114 10616 16120 10628
rect 16172 10616 16178 10668
rect 16758 10616 16764 10668
rect 16816 10616 16822 10668
rect 17494 10616 17500 10668
rect 17552 10656 17558 10668
rect 17865 10659 17923 10665
rect 17865 10656 17877 10659
rect 17552 10628 17877 10656
rect 17552 10616 17558 10628
rect 17865 10625 17877 10628
rect 17911 10625 17923 10659
rect 17865 10619 17923 10625
rect 19150 10616 19156 10668
rect 19208 10656 19214 10668
rect 21008 10665 21036 10764
rect 22554 10752 22560 10764
rect 22612 10752 22618 10804
rect 22278 10684 22284 10736
rect 22336 10684 22342 10736
rect 22738 10684 22744 10736
rect 22796 10684 22802 10736
rect 20993 10659 21051 10665
rect 19208 10628 19274 10656
rect 19208 10616 19214 10628
rect 20993 10625 21005 10659
rect 21039 10625 21051 10659
rect 20993 10619 21051 10625
rect 21174 10616 21180 10668
rect 21232 10656 21238 10668
rect 21726 10656 21732 10668
rect 21232 10628 21732 10656
rect 21232 10616 21238 10628
rect 21726 10616 21732 10628
rect 21784 10616 21790 10668
rect 11103 10560 12112 10588
rect 12253 10591 12311 10597
rect 11103 10557 11115 10560
rect 11057 10551 11115 10557
rect 12253 10557 12265 10591
rect 12299 10557 12311 10591
rect 12253 10551 12311 10557
rect 14093 10591 14151 10597
rect 14093 10557 14105 10591
rect 14139 10557 14151 10591
rect 14093 10551 14151 10557
rect 14185 10591 14243 10597
rect 14185 10557 14197 10591
rect 14231 10557 14243 10591
rect 14185 10551 14243 10557
rect 15381 10591 15439 10597
rect 15381 10557 15393 10591
rect 15427 10557 15439 10591
rect 15381 10551 15439 10557
rect 18141 10591 18199 10597
rect 18141 10557 18153 10591
rect 18187 10588 18199 10591
rect 18782 10588 18788 10600
rect 18187 10560 18788 10588
rect 18187 10557 18199 10560
rect 18141 10551 18199 10557
rect 6546 10520 6552 10532
rect 5092 10492 6552 10520
rect 4801 10483 4859 10489
rect 2498 10412 2504 10464
rect 2556 10452 2562 10464
rect 2593 10455 2651 10461
rect 2593 10452 2605 10455
rect 2556 10424 2605 10452
rect 2556 10412 2562 10424
rect 2593 10421 2605 10424
rect 2639 10421 2651 10455
rect 4816 10452 4844 10483
rect 6546 10480 6552 10492
rect 6604 10480 6610 10532
rect 9490 10480 9496 10532
rect 9548 10520 9554 10532
rect 9585 10523 9643 10529
rect 9585 10520 9597 10523
rect 9548 10492 9597 10520
rect 9548 10480 9554 10492
rect 9585 10489 9597 10492
rect 9631 10520 9643 10523
rect 12158 10520 12164 10532
rect 9631 10492 12164 10520
rect 9631 10489 9643 10492
rect 9585 10483 9643 10489
rect 12158 10480 12164 10492
rect 12216 10480 12222 10532
rect 14108 10520 14136 10551
rect 12268 10492 14136 10520
rect 14200 10520 14228 10551
rect 15396 10520 15424 10551
rect 18782 10548 18788 10560
rect 18840 10548 18846 10600
rect 19610 10548 19616 10600
rect 19668 10588 19674 10600
rect 22005 10591 22063 10597
rect 22005 10588 22017 10591
rect 19668 10560 22017 10588
rect 19668 10548 19674 10560
rect 22005 10557 22017 10560
rect 22051 10557 22063 10591
rect 22005 10551 22063 10557
rect 16022 10520 16028 10532
rect 14200 10492 16028 10520
rect 4890 10452 4896 10464
rect 4816 10424 4896 10452
rect 2593 10415 2651 10421
rect 4890 10412 4896 10424
rect 4948 10452 4954 10464
rect 5442 10452 5448 10464
rect 4948 10424 5448 10452
rect 4948 10412 4954 10424
rect 5442 10412 5448 10424
rect 5500 10412 5506 10464
rect 5626 10412 5632 10464
rect 5684 10412 5690 10464
rect 5718 10412 5724 10464
rect 5776 10452 5782 10464
rect 6362 10452 6368 10464
rect 5776 10424 6368 10452
rect 5776 10412 5782 10424
rect 6362 10412 6368 10424
rect 6420 10452 6426 10464
rect 6641 10455 6699 10461
rect 6641 10452 6653 10455
rect 6420 10424 6653 10452
rect 6420 10412 6426 10424
rect 6641 10421 6653 10424
rect 6687 10421 6699 10455
rect 6641 10415 6699 10421
rect 9398 10412 9404 10464
rect 9456 10452 9462 10464
rect 10778 10452 10784 10464
rect 9456 10424 10784 10452
rect 9456 10412 9462 10424
rect 10778 10412 10784 10424
rect 10836 10412 10842 10464
rect 11146 10412 11152 10464
rect 11204 10452 11210 10464
rect 12268 10452 12296 10492
rect 11204 10424 12296 10452
rect 11204 10412 11210 10424
rect 12342 10412 12348 10464
rect 12400 10452 12406 10464
rect 14200 10452 14228 10492
rect 15212 10464 15240 10492
rect 16022 10480 16028 10492
rect 16080 10480 16086 10532
rect 12400 10424 14228 10452
rect 12400 10412 12406 10424
rect 14458 10412 14464 10464
rect 14516 10452 14522 10464
rect 14645 10455 14703 10461
rect 14645 10452 14657 10455
rect 14516 10424 14657 10452
rect 14516 10412 14522 10424
rect 14645 10421 14657 10424
rect 14691 10421 14703 10455
rect 14645 10415 14703 10421
rect 15194 10412 15200 10464
rect 15252 10412 15258 10464
rect 16942 10412 16948 10464
rect 17000 10412 17006 10464
rect 18690 10412 18696 10464
rect 18748 10452 18754 10464
rect 19613 10455 19671 10461
rect 19613 10452 19625 10455
rect 18748 10424 19625 10452
rect 18748 10412 18754 10424
rect 19613 10421 19625 10424
rect 19659 10421 19671 10455
rect 19613 10415 19671 10421
rect 21174 10412 21180 10464
rect 21232 10412 21238 10464
rect 23753 10455 23811 10461
rect 23753 10421 23765 10455
rect 23799 10452 23811 10455
rect 23842 10452 23848 10464
rect 23799 10424 23848 10452
rect 23799 10421 23811 10424
rect 23753 10415 23811 10421
rect 23842 10412 23848 10424
rect 23900 10412 23906 10464
rect 1104 10362 25852 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 12214 10362
rect 12266 10310 12278 10362
rect 12330 10310 12342 10362
rect 12394 10310 12406 10362
rect 12458 10310 12470 10362
rect 12522 10310 20214 10362
rect 20266 10310 20278 10362
rect 20330 10310 20342 10362
rect 20394 10310 20406 10362
rect 20458 10310 20470 10362
rect 20522 10310 25852 10362
rect 1104 10288 25852 10310
rect 5445 10251 5503 10257
rect 5445 10217 5457 10251
rect 5491 10248 5503 10251
rect 6454 10248 6460 10260
rect 5491 10220 6460 10248
rect 5491 10217 5503 10220
rect 5445 10211 5503 10217
rect 6454 10208 6460 10220
rect 6512 10208 6518 10260
rect 6914 10208 6920 10260
rect 6972 10208 6978 10260
rect 7926 10208 7932 10260
rect 7984 10208 7990 10260
rect 9030 10208 9036 10260
rect 9088 10208 9094 10260
rect 9214 10208 9220 10260
rect 9272 10248 9278 10260
rect 9272 10220 12434 10248
rect 9272 10208 9278 10220
rect 3970 10140 3976 10192
rect 4028 10180 4034 10192
rect 4157 10183 4215 10189
rect 4157 10180 4169 10183
rect 4028 10152 4169 10180
rect 4028 10140 4034 10152
rect 4157 10149 4169 10152
rect 4203 10180 4215 10183
rect 5718 10180 5724 10192
rect 4203 10152 4752 10180
rect 4203 10149 4215 10152
rect 4157 10143 4215 10149
rect 4246 10072 4252 10124
rect 4304 10112 4310 10124
rect 4617 10115 4675 10121
rect 4617 10112 4629 10115
rect 4304 10084 4629 10112
rect 4304 10072 4310 10084
rect 4617 10081 4629 10084
rect 4663 10081 4675 10115
rect 4617 10075 4675 10081
rect 1486 10004 1492 10056
rect 1544 10004 1550 10056
rect 1762 9936 1768 9988
rect 1820 9936 1826 9988
rect 2498 9936 2504 9988
rect 2556 9936 2562 9988
rect 3881 9979 3939 9985
rect 3881 9945 3893 9979
rect 3927 9976 3939 9979
rect 4154 9976 4160 9988
rect 3927 9948 4160 9976
rect 3927 9945 3939 9948
rect 3881 9939 3939 9945
rect 4154 9936 4160 9948
rect 4212 9976 4218 9988
rect 4430 9976 4436 9988
rect 4212 9948 4436 9976
rect 4212 9936 4218 9948
rect 4430 9936 4436 9948
rect 4488 9936 4494 9988
rect 4724 9976 4752 10152
rect 4908 10152 5724 10180
rect 4908 10121 4936 10152
rect 5718 10140 5724 10152
rect 5776 10140 5782 10192
rect 7561 10183 7619 10189
rect 7561 10180 7573 10183
rect 6104 10152 7573 10180
rect 6104 10124 6132 10152
rect 7561 10149 7573 10152
rect 7607 10149 7619 10183
rect 10318 10180 10324 10192
rect 7561 10143 7619 10149
rect 8588 10152 10324 10180
rect 4893 10115 4951 10121
rect 4893 10081 4905 10115
rect 4939 10081 4951 10115
rect 6086 10112 6092 10124
rect 4893 10075 4951 10081
rect 5000 10084 6092 10112
rect 5000 10053 5028 10084
rect 6086 10072 6092 10084
rect 6144 10072 6150 10124
rect 6454 10072 6460 10124
rect 6512 10112 6518 10124
rect 8588 10121 8616 10152
rect 9692 10124 9720 10152
rect 10318 10140 10324 10152
rect 10376 10140 10382 10192
rect 12406 10180 12434 10220
rect 12618 10208 12624 10260
rect 12676 10208 12682 10260
rect 14918 10208 14924 10260
rect 14976 10208 14982 10260
rect 16758 10208 16764 10260
rect 16816 10248 16822 10260
rect 16945 10251 17003 10257
rect 16945 10248 16957 10251
rect 16816 10220 16957 10248
rect 16816 10208 16822 10220
rect 16945 10217 16957 10220
rect 16991 10217 17003 10251
rect 16945 10211 17003 10217
rect 19150 10208 19156 10260
rect 19208 10248 19214 10260
rect 19337 10251 19395 10257
rect 19337 10248 19349 10251
rect 19208 10220 19349 10248
rect 19208 10208 19214 10220
rect 19337 10217 19349 10220
rect 19383 10217 19395 10251
rect 19337 10211 19395 10217
rect 22738 10208 22744 10260
rect 22796 10208 22802 10260
rect 15286 10180 15292 10192
rect 12406 10152 15292 10180
rect 15286 10140 15292 10152
rect 15344 10140 15350 10192
rect 16209 10183 16267 10189
rect 16209 10180 16221 10183
rect 15580 10152 16221 10180
rect 8573 10115 8631 10121
rect 6512 10084 7512 10112
rect 6512 10072 6518 10084
rect 4985 10047 5043 10053
rect 4985 10013 4997 10047
rect 5031 10013 5043 10047
rect 4985 10007 5043 10013
rect 5442 10004 5448 10056
rect 5500 10044 5506 10056
rect 5629 10047 5687 10053
rect 5629 10044 5641 10047
rect 5500 10016 5641 10044
rect 5500 10004 5506 10016
rect 5629 10013 5641 10016
rect 5675 10044 5687 10047
rect 5810 10044 5816 10056
rect 5675 10016 5816 10044
rect 5675 10013 5687 10016
rect 5629 10007 5687 10013
rect 5810 10004 5816 10016
rect 5868 10004 5874 10056
rect 5902 10004 5908 10056
rect 5960 10004 5966 10056
rect 6178 10004 6184 10056
rect 6236 10004 6242 10056
rect 6270 10004 6276 10056
rect 6328 10044 6334 10056
rect 6549 10047 6607 10053
rect 6328 10016 6373 10044
rect 6328 10004 6334 10016
rect 6549 10013 6561 10047
rect 6595 10044 6607 10047
rect 6825 10047 6883 10053
rect 6825 10044 6837 10047
rect 6595 10016 6837 10044
rect 6595 10013 6607 10016
rect 6549 10007 6607 10013
rect 6825 10013 6837 10016
rect 6871 10013 6883 10047
rect 6825 10007 6883 10013
rect 6914 10004 6920 10056
rect 6972 10044 6978 10056
rect 7484 10053 7512 10084
rect 8573 10081 8585 10115
rect 8619 10081 8631 10115
rect 8573 10075 8631 10081
rect 9490 10072 9496 10124
rect 9548 10072 9554 10124
rect 9674 10072 9680 10124
rect 9732 10112 9738 10124
rect 9732 10084 9757 10112
rect 9732 10072 9738 10084
rect 10410 10072 10416 10124
rect 10468 10072 10474 10124
rect 11238 10072 11244 10124
rect 11296 10112 11302 10124
rect 12894 10112 12900 10124
rect 11296 10084 12480 10112
rect 11296 10072 11302 10084
rect 7193 10047 7251 10053
rect 7193 10044 7205 10047
rect 6972 10016 7205 10044
rect 6972 10004 6978 10016
rect 7193 10013 7205 10016
rect 7239 10013 7251 10047
rect 7193 10007 7251 10013
rect 7469 10047 7527 10053
rect 7469 10013 7481 10047
rect 7515 10013 7527 10047
rect 7469 10007 7527 10013
rect 7558 10004 7564 10056
rect 7616 10044 7622 10056
rect 7653 10047 7711 10053
rect 7653 10044 7665 10047
rect 7616 10016 7665 10044
rect 7616 10004 7622 10016
rect 7653 10013 7665 10016
rect 7699 10013 7711 10047
rect 7653 10007 7711 10013
rect 7926 10004 7932 10056
rect 7984 10044 7990 10056
rect 12452 10053 12480 10084
rect 12636 10084 12900 10112
rect 12636 10053 12664 10084
rect 12894 10072 12900 10084
rect 12952 10072 12958 10124
rect 15102 10072 15108 10124
rect 15160 10112 15166 10124
rect 15580 10121 15608 10152
rect 16209 10149 16221 10152
rect 16255 10180 16267 10183
rect 16255 10152 17632 10180
rect 16255 10149 16267 10152
rect 16209 10143 16267 10149
rect 15381 10115 15439 10121
rect 15381 10112 15393 10115
rect 15160 10084 15393 10112
rect 15160 10072 15166 10084
rect 15381 10081 15393 10084
rect 15427 10081 15439 10115
rect 15381 10075 15439 10081
rect 15565 10115 15623 10121
rect 15565 10081 15577 10115
rect 15611 10081 15623 10115
rect 15565 10075 15623 10081
rect 16574 10072 16580 10124
rect 16632 10112 16638 10124
rect 17604 10121 17632 10152
rect 19352 10152 20300 10180
rect 17405 10115 17463 10121
rect 17405 10112 17417 10115
rect 16632 10084 17417 10112
rect 16632 10072 16638 10084
rect 17405 10081 17417 10084
rect 17451 10081 17463 10115
rect 17405 10075 17463 10081
rect 17589 10115 17647 10121
rect 17589 10081 17601 10115
rect 17635 10112 17647 10115
rect 18230 10112 18236 10124
rect 17635 10084 18236 10112
rect 17635 10081 17647 10084
rect 17589 10075 17647 10081
rect 18230 10072 18236 10084
rect 18288 10072 18294 10124
rect 9401 10047 9459 10053
rect 9401 10044 9413 10047
rect 7984 10016 9413 10044
rect 7984 10004 7990 10016
rect 9401 10013 9413 10016
rect 9447 10013 9459 10047
rect 9401 10007 9459 10013
rect 12437 10047 12495 10053
rect 12437 10013 12449 10047
rect 12483 10013 12495 10047
rect 12437 10007 12495 10013
rect 12621 10047 12679 10053
rect 12621 10013 12633 10047
rect 12667 10013 12679 10047
rect 12621 10007 12679 10013
rect 5534 9976 5540 9988
rect 4724 9948 5540 9976
rect 5534 9936 5540 9948
rect 5592 9936 5598 9988
rect 6086 9936 6092 9988
rect 6144 9976 6150 9988
rect 8297 9979 8355 9985
rect 6144 9948 7052 9976
rect 6144 9936 6150 9948
rect 3234 9868 3240 9920
rect 3292 9868 3298 9920
rect 4341 9911 4399 9917
rect 4341 9877 4353 9911
rect 4387 9908 4399 9911
rect 5350 9908 5356 9920
rect 4387 9880 5356 9908
rect 4387 9877 4399 9880
rect 4341 9871 4399 9877
rect 5350 9868 5356 9880
rect 5408 9868 5414 9920
rect 5813 9911 5871 9917
rect 5813 9877 5825 9911
rect 5859 9908 5871 9911
rect 6546 9908 6552 9920
rect 5859 9880 6552 9908
rect 5859 9877 5871 9880
rect 5813 9871 5871 9877
rect 6546 9868 6552 9880
rect 6604 9868 6610 9920
rect 6638 9868 6644 9920
rect 6696 9908 6702 9920
rect 7024 9917 7052 9948
rect 8297 9945 8309 9979
rect 8343 9976 8355 9979
rect 8754 9976 8760 9988
rect 8343 9948 8760 9976
rect 8343 9945 8355 9948
rect 8297 9939 8355 9945
rect 8754 9936 8760 9948
rect 8812 9936 8818 9988
rect 10686 9936 10692 9988
rect 10744 9936 10750 9988
rect 11974 9976 11980 9988
rect 11914 9948 11980 9976
rect 11974 9936 11980 9948
rect 12032 9936 12038 9988
rect 12636 9976 12664 10007
rect 12710 10004 12716 10056
rect 12768 10044 12774 10056
rect 13357 10047 13415 10053
rect 13357 10044 13369 10047
rect 12768 10016 13369 10044
rect 12768 10004 12774 10016
rect 13357 10013 13369 10016
rect 13403 10044 13415 10047
rect 14277 10047 14335 10053
rect 14277 10044 14289 10047
rect 13403 10016 14289 10044
rect 13403 10013 13415 10016
rect 13357 10007 13415 10013
rect 14277 10013 14289 10016
rect 14323 10013 14335 10047
rect 14277 10007 14335 10013
rect 14384 10016 15516 10044
rect 14384 9976 14412 10016
rect 12084 9948 12664 9976
rect 13188 9948 14412 9976
rect 14461 9979 14519 9985
rect 6917 9911 6975 9917
rect 6917 9908 6929 9911
rect 6696 9880 6929 9908
rect 6696 9868 6702 9880
rect 6917 9877 6929 9880
rect 6963 9877 6975 9911
rect 6917 9871 6975 9877
rect 7009 9911 7067 9917
rect 7009 9877 7021 9911
rect 7055 9877 7067 9911
rect 7009 9871 7067 9877
rect 8389 9911 8447 9917
rect 8389 9877 8401 9911
rect 8435 9908 8447 9911
rect 9214 9908 9220 9920
rect 8435 9880 9220 9908
rect 8435 9877 8447 9880
rect 8389 9871 8447 9877
rect 9214 9868 9220 9880
rect 9272 9868 9278 9920
rect 11698 9868 11704 9920
rect 11756 9908 11762 9920
rect 12084 9908 12112 9948
rect 11756 9880 12112 9908
rect 11756 9868 11762 9880
rect 12158 9868 12164 9920
rect 12216 9868 12222 9920
rect 13078 9868 13084 9920
rect 13136 9908 13142 9920
rect 13188 9917 13216 9948
rect 14461 9945 14473 9979
rect 14507 9976 14519 9979
rect 15378 9976 15384 9988
rect 14507 9948 15384 9976
rect 14507 9945 14519 9948
rect 14461 9939 14519 9945
rect 15378 9936 15384 9948
rect 15436 9936 15442 9988
rect 13173 9911 13231 9917
rect 13173 9908 13185 9911
rect 13136 9880 13185 9908
rect 13136 9868 13142 9880
rect 13173 9877 13185 9880
rect 13219 9877 13231 9911
rect 13173 9871 13231 9877
rect 15286 9868 15292 9920
rect 15344 9868 15350 9920
rect 15488 9908 15516 10016
rect 16022 10004 16028 10056
rect 16080 10004 16086 10056
rect 16114 10004 16120 10056
rect 16172 10044 16178 10056
rect 18325 10047 18383 10053
rect 18325 10044 18337 10047
rect 16172 10016 18337 10044
rect 16172 10004 16178 10016
rect 18325 10013 18337 10016
rect 18371 10013 18383 10047
rect 18325 10007 18383 10013
rect 18417 10047 18475 10053
rect 18417 10013 18429 10047
rect 18463 10044 18475 10047
rect 18690 10044 18696 10056
rect 18463 10016 18696 10044
rect 18463 10013 18475 10016
rect 18417 10007 18475 10013
rect 18690 10004 18696 10016
rect 18748 10004 18754 10056
rect 19150 10004 19156 10056
rect 19208 10044 19214 10056
rect 19352 10053 19380 10152
rect 19610 10072 19616 10124
rect 19668 10112 19674 10124
rect 20165 10115 20223 10121
rect 20165 10112 20177 10115
rect 19668 10084 20177 10112
rect 19668 10072 19674 10084
rect 20165 10081 20177 10084
rect 20211 10081 20223 10115
rect 20272 10112 20300 10152
rect 23382 10140 23388 10192
rect 23440 10180 23446 10192
rect 23440 10152 23612 10180
rect 23440 10140 23446 10152
rect 21082 10112 21088 10124
rect 20272 10084 21088 10112
rect 20165 10075 20223 10081
rect 21082 10072 21088 10084
rect 21140 10072 21146 10124
rect 21450 10072 21456 10124
rect 21508 10112 21514 10124
rect 23584 10121 23612 10152
rect 23477 10115 23535 10121
rect 23477 10112 23489 10115
rect 21508 10084 23489 10112
rect 21508 10072 21514 10084
rect 23477 10081 23489 10084
rect 23523 10081 23535 10115
rect 23477 10075 23535 10081
rect 23569 10115 23627 10121
rect 23569 10081 23581 10115
rect 23615 10081 23627 10115
rect 23569 10075 23627 10081
rect 19337 10047 19395 10053
rect 19337 10044 19349 10047
rect 19208 10016 19349 10044
rect 19208 10004 19214 10016
rect 19337 10013 19349 10016
rect 19383 10013 19395 10047
rect 19337 10007 19395 10013
rect 19518 10004 19524 10056
rect 19576 10004 19582 10056
rect 22554 10004 22560 10056
rect 22612 10004 22618 10056
rect 22741 10047 22799 10053
rect 22741 10013 22753 10047
rect 22787 10044 22799 10047
rect 24118 10044 24124 10056
rect 22787 10016 24124 10044
rect 22787 10013 22799 10016
rect 22741 10007 22799 10013
rect 17313 9979 17371 9985
rect 17313 9945 17325 9979
rect 17359 9976 17371 9979
rect 17770 9976 17776 9988
rect 17359 9948 17776 9976
rect 17359 9945 17371 9948
rect 17313 9939 17371 9945
rect 17770 9936 17776 9948
rect 17828 9936 17834 9988
rect 18708 9948 19380 9976
rect 18708 9908 18736 9948
rect 15488 9880 18736 9908
rect 18785 9911 18843 9917
rect 18785 9877 18797 9911
rect 18831 9908 18843 9911
rect 18966 9908 18972 9920
rect 18831 9880 18972 9908
rect 18831 9877 18843 9880
rect 18785 9871 18843 9877
rect 18966 9868 18972 9880
rect 19024 9868 19030 9920
rect 19352 9908 19380 9948
rect 20070 9936 20076 9988
rect 20128 9976 20134 9988
rect 20441 9979 20499 9985
rect 20441 9976 20453 9979
rect 20128 9948 20453 9976
rect 20128 9936 20134 9948
rect 20441 9945 20453 9948
rect 20487 9945 20499 9979
rect 20441 9939 20499 9945
rect 21174 9936 21180 9988
rect 21232 9936 21238 9988
rect 22756 9976 22784 10007
rect 24118 10004 24124 10016
rect 24176 10004 24182 10056
rect 21836 9948 22784 9976
rect 23385 9979 23443 9985
rect 21836 9908 21864 9948
rect 23385 9945 23397 9979
rect 23431 9976 23443 9979
rect 24762 9976 24768 9988
rect 23431 9948 24768 9976
rect 23431 9945 23443 9948
rect 23385 9939 23443 9945
rect 24762 9936 24768 9948
rect 24820 9936 24826 9988
rect 19352 9880 21864 9908
rect 21910 9868 21916 9920
rect 21968 9868 21974 9920
rect 22738 9868 22744 9920
rect 22796 9908 22802 9920
rect 23017 9911 23075 9917
rect 23017 9908 23029 9911
rect 22796 9880 23029 9908
rect 22796 9868 22802 9880
rect 23017 9877 23029 9880
rect 23063 9877 23075 9911
rect 23017 9871 23075 9877
rect 1104 9818 25852 9840
rect 1104 9766 8214 9818
rect 8266 9766 8278 9818
rect 8330 9766 8342 9818
rect 8394 9766 8406 9818
rect 8458 9766 8470 9818
rect 8522 9766 16214 9818
rect 16266 9766 16278 9818
rect 16330 9766 16342 9818
rect 16394 9766 16406 9818
rect 16458 9766 16470 9818
rect 16522 9766 24214 9818
rect 24266 9766 24278 9818
rect 24330 9766 24342 9818
rect 24394 9766 24406 9818
rect 24458 9766 24470 9818
rect 24522 9766 25852 9818
rect 1104 9744 25852 9766
rect 1762 9664 1768 9716
rect 1820 9704 1826 9716
rect 2041 9707 2099 9713
rect 2041 9704 2053 9707
rect 1820 9676 2053 9704
rect 1820 9664 1826 9676
rect 2041 9673 2053 9676
rect 2087 9673 2099 9707
rect 2041 9667 2099 9673
rect 2961 9707 3019 9713
rect 2961 9673 2973 9707
rect 3007 9704 3019 9707
rect 3234 9704 3240 9716
rect 3007 9676 3240 9704
rect 3007 9673 3019 9676
rect 2961 9667 3019 9673
rect 3234 9664 3240 9676
rect 3292 9664 3298 9716
rect 5902 9664 5908 9716
rect 5960 9704 5966 9716
rect 5960 9676 6776 9704
rect 5960 9664 5966 9676
rect 3053 9639 3111 9645
rect 3053 9605 3065 9639
rect 3099 9636 3111 9639
rect 4246 9636 4252 9648
rect 3099 9608 4252 9636
rect 3099 9605 3111 9608
rect 3053 9599 3111 9605
rect 4246 9596 4252 9608
rect 4304 9596 4310 9648
rect 4430 9596 4436 9648
rect 4488 9636 4494 9648
rect 4488 9608 5856 9636
rect 4488 9596 4494 9608
rect 2225 9571 2283 9577
rect 2225 9537 2237 9571
rect 2271 9568 2283 9571
rect 4341 9571 4399 9577
rect 2271 9540 2636 9568
rect 2271 9537 2283 9540
rect 2225 9531 2283 9537
rect 2608 9441 2636 9540
rect 4341 9537 4353 9571
rect 4387 9568 4399 9571
rect 4522 9568 4528 9580
rect 4387 9540 4528 9568
rect 4387 9537 4399 9540
rect 4341 9531 4399 9537
rect 4522 9528 4528 9540
rect 4580 9528 4586 9580
rect 4617 9571 4675 9577
rect 4617 9537 4629 9571
rect 4663 9568 4675 9571
rect 4985 9571 5043 9577
rect 4985 9568 4997 9571
rect 4663 9540 4997 9568
rect 4663 9537 4675 9540
rect 4617 9531 4675 9537
rect 4985 9537 4997 9540
rect 5031 9537 5043 9571
rect 4985 9531 5043 9537
rect 5169 9571 5227 9577
rect 5169 9537 5181 9571
rect 5215 9568 5227 9571
rect 5215 9540 5304 9568
rect 5215 9537 5227 9540
rect 5169 9531 5227 9537
rect 3237 9503 3295 9509
rect 3237 9469 3249 9503
rect 3283 9500 3295 9503
rect 3418 9500 3424 9512
rect 3283 9472 3424 9500
rect 3283 9469 3295 9472
rect 3237 9463 3295 9469
rect 3418 9460 3424 9472
rect 3476 9460 3482 9512
rect 2593 9435 2651 9441
rect 2593 9401 2605 9435
rect 2639 9401 2651 9435
rect 2593 9395 2651 9401
rect 3970 9392 3976 9444
rect 4028 9432 4034 9444
rect 4433 9435 4491 9441
rect 4433 9432 4445 9435
rect 4028 9404 4445 9432
rect 4028 9392 4034 9404
rect 4433 9401 4445 9404
rect 4479 9401 4491 9435
rect 4433 9395 4491 9401
rect 4525 9435 4583 9441
rect 4525 9401 4537 9435
rect 4571 9432 4583 9435
rect 4706 9432 4712 9444
rect 4571 9404 4712 9432
rect 4571 9401 4583 9404
rect 4525 9395 4583 9401
rect 4706 9392 4712 9404
rect 4764 9432 4770 9444
rect 4982 9432 4988 9444
rect 4764 9404 4988 9432
rect 4764 9392 4770 9404
rect 4982 9392 4988 9404
rect 5040 9392 5046 9444
rect 4062 9324 4068 9376
rect 4120 9364 4126 9376
rect 4157 9367 4215 9373
rect 4157 9364 4169 9367
rect 4120 9336 4169 9364
rect 4120 9324 4126 9336
rect 4157 9333 4169 9336
rect 4203 9333 4215 9367
rect 5276 9364 5304 9540
rect 5350 9528 5356 9580
rect 5408 9528 5414 9580
rect 5445 9571 5503 9577
rect 5445 9537 5457 9571
rect 5491 9568 5503 9571
rect 5626 9568 5632 9580
rect 5491 9540 5632 9568
rect 5491 9537 5503 9540
rect 5445 9531 5503 9537
rect 5626 9528 5632 9540
rect 5684 9528 5690 9580
rect 5718 9528 5724 9580
rect 5776 9528 5782 9580
rect 5828 9577 5856 9608
rect 6086 9596 6092 9648
rect 6144 9596 6150 9648
rect 6546 9596 6552 9648
rect 6604 9596 6610 9648
rect 6748 9580 6776 9676
rect 9214 9664 9220 9716
rect 9272 9664 9278 9716
rect 10229 9707 10287 9713
rect 10229 9673 10241 9707
rect 10275 9704 10287 9707
rect 10686 9704 10692 9716
rect 10275 9676 10692 9704
rect 10275 9673 10287 9676
rect 10229 9667 10287 9673
rect 10686 9664 10692 9676
rect 10744 9664 10750 9716
rect 15286 9664 15292 9716
rect 15344 9704 15350 9716
rect 15933 9707 15991 9713
rect 15933 9704 15945 9707
rect 15344 9676 15945 9704
rect 15344 9664 15350 9676
rect 15933 9673 15945 9676
rect 15979 9673 15991 9707
rect 15933 9667 15991 9673
rect 18782 9664 18788 9716
rect 18840 9664 18846 9716
rect 19518 9664 19524 9716
rect 19576 9704 19582 9716
rect 19576 9676 22048 9704
rect 19576 9664 19582 9676
rect 7834 9636 7840 9648
rect 7484 9608 7840 9636
rect 5814 9571 5872 9577
rect 5814 9537 5826 9571
rect 5860 9537 5872 9571
rect 5814 9531 5872 9537
rect 5902 9528 5908 9580
rect 5960 9568 5966 9580
rect 6270 9568 6276 9580
rect 5960 9540 6276 9568
rect 5960 9528 5966 9540
rect 6270 9528 6276 9540
rect 6328 9568 6334 9580
rect 6457 9571 6515 9577
rect 6457 9568 6469 9571
rect 6328 9540 6469 9568
rect 6328 9528 6334 9540
rect 6457 9537 6469 9540
rect 6503 9537 6515 9571
rect 6457 9531 6515 9537
rect 6730 9528 6736 9580
rect 6788 9528 6794 9580
rect 7190 9528 7196 9580
rect 7248 9568 7254 9580
rect 7484 9577 7512 9608
rect 7834 9596 7840 9608
rect 7892 9596 7898 9648
rect 9306 9636 9312 9648
rect 8970 9608 9312 9636
rect 9306 9596 9312 9608
rect 9364 9596 9370 9648
rect 9858 9596 9864 9648
rect 9916 9636 9922 9648
rect 10778 9636 10784 9648
rect 9916 9608 10784 9636
rect 9916 9596 9922 9608
rect 10778 9596 10784 9608
rect 10836 9636 10842 9648
rect 11698 9636 11704 9648
rect 10836 9608 11704 9636
rect 10836 9596 10842 9608
rect 7469 9571 7527 9577
rect 7469 9568 7481 9571
rect 7248 9540 7481 9568
rect 7248 9528 7254 9540
rect 7469 9537 7481 9540
rect 7515 9537 7527 9571
rect 7469 9531 7527 9537
rect 10045 9571 10103 9577
rect 10045 9537 10057 9571
rect 10091 9568 10103 9571
rect 10410 9568 10416 9580
rect 10091 9540 10416 9568
rect 10091 9537 10103 9540
rect 10045 9531 10103 9537
rect 10410 9528 10416 9540
rect 10468 9528 10474 9580
rect 10686 9528 10692 9580
rect 10744 9528 10750 9580
rect 11072 9577 11100 9608
rect 11698 9596 11704 9608
rect 11756 9636 11762 9648
rect 11756 9608 11928 9636
rect 11756 9596 11762 9608
rect 11057 9571 11115 9577
rect 11057 9537 11069 9571
rect 11103 9537 11115 9571
rect 11057 9531 11115 9537
rect 11238 9528 11244 9580
rect 11296 9528 11302 9580
rect 11900 9577 11928 9608
rect 11974 9596 11980 9648
rect 12032 9596 12038 9648
rect 14458 9596 14464 9648
rect 14516 9596 14522 9648
rect 15470 9596 15476 9648
rect 15528 9596 15534 9648
rect 16942 9596 16948 9648
rect 17000 9636 17006 9648
rect 17037 9639 17095 9645
rect 17037 9636 17049 9639
rect 17000 9608 17049 9636
rect 17000 9596 17006 9608
rect 17037 9605 17049 9608
rect 17083 9605 17095 9639
rect 17037 9599 17095 9605
rect 17678 9596 17684 9648
rect 17736 9596 17742 9648
rect 22020 9636 22048 9676
rect 22554 9664 22560 9716
rect 22612 9704 22618 9716
rect 23474 9704 23480 9716
rect 22612 9676 23480 9704
rect 22612 9664 22618 9676
rect 23474 9664 23480 9676
rect 23532 9664 23538 9716
rect 22020 9608 23060 9636
rect 23032 9580 23060 9608
rect 11885 9571 11943 9577
rect 11885 9537 11897 9571
rect 11931 9537 11943 9571
rect 11885 9531 11943 9537
rect 12066 9528 12072 9580
rect 12124 9528 12130 9580
rect 18966 9528 18972 9580
rect 19024 9528 19030 9580
rect 19518 9528 19524 9580
rect 19576 9528 19582 9580
rect 20898 9528 20904 9580
rect 20956 9528 20962 9580
rect 22094 9528 22100 9580
rect 22152 9528 22158 9580
rect 22557 9571 22615 9577
rect 22557 9537 22569 9571
rect 22603 9568 22615 9571
rect 22738 9568 22744 9580
rect 22603 9540 22744 9568
rect 22603 9537 22615 9540
rect 22557 9531 22615 9537
rect 22738 9528 22744 9540
rect 22796 9528 22802 9580
rect 23014 9528 23020 9580
rect 23072 9528 23078 9580
rect 24394 9528 24400 9580
rect 24452 9528 24458 9580
rect 5644 9500 5672 9528
rect 6822 9500 6828 9512
rect 5644 9472 6828 9500
rect 6822 9460 6828 9472
rect 6880 9460 6886 9512
rect 7742 9460 7748 9512
rect 7800 9460 7806 9512
rect 13170 9460 13176 9512
rect 13228 9500 13234 9512
rect 14185 9503 14243 9509
rect 14185 9500 14197 9503
rect 13228 9472 14197 9500
rect 13228 9460 13234 9472
rect 14185 9469 14197 9472
rect 14231 9469 14243 9503
rect 14185 9463 14243 9469
rect 16666 9460 16672 9512
rect 16724 9500 16730 9512
rect 16761 9503 16819 9509
rect 16761 9500 16773 9503
rect 16724 9472 16773 9500
rect 16724 9460 16730 9472
rect 16761 9469 16773 9472
rect 16807 9469 16819 9503
rect 16761 9463 16819 9469
rect 17770 9460 17776 9512
rect 17828 9500 17834 9512
rect 18509 9503 18567 9509
rect 18509 9500 18521 9503
rect 17828 9472 18521 9500
rect 17828 9460 17834 9472
rect 18509 9469 18521 9472
rect 18555 9469 18567 9503
rect 18509 9463 18567 9469
rect 19794 9460 19800 9512
rect 19852 9460 19858 9512
rect 21269 9503 21327 9509
rect 21269 9469 21281 9503
rect 21315 9500 21327 9503
rect 21450 9500 21456 9512
rect 21315 9472 21456 9500
rect 21315 9469 21327 9472
rect 21269 9463 21327 9469
rect 21450 9460 21456 9472
rect 21508 9460 21514 9512
rect 23293 9503 23351 9509
rect 23293 9500 23305 9503
rect 22756 9472 23305 9500
rect 11054 9392 11060 9444
rect 11112 9392 11118 9444
rect 22756 9441 22784 9472
rect 23293 9469 23305 9472
rect 23339 9469 23351 9503
rect 23293 9463 23351 9469
rect 24762 9460 24768 9512
rect 24820 9460 24826 9512
rect 22741 9435 22799 9441
rect 22741 9401 22753 9435
rect 22787 9401 22799 9435
rect 22741 9395 22799 9401
rect 5905 9367 5963 9373
rect 5905 9364 5917 9367
rect 5276 9336 5917 9364
rect 4157 9327 4215 9333
rect 5905 9333 5917 9336
rect 5951 9333 5963 9367
rect 5905 9327 5963 9333
rect 6641 9367 6699 9373
rect 6641 9333 6653 9367
rect 6687 9364 6699 9367
rect 7558 9364 7564 9376
rect 6687 9336 7564 9364
rect 6687 9333 6699 9336
rect 6641 9327 6699 9333
rect 7558 9324 7564 9336
rect 7616 9324 7622 9376
rect 9582 9324 9588 9376
rect 9640 9364 9646 9376
rect 10505 9367 10563 9373
rect 10505 9364 10517 9367
rect 9640 9336 10517 9364
rect 9640 9324 9646 9336
rect 10505 9333 10517 9336
rect 10551 9333 10563 9367
rect 10505 9327 10563 9333
rect 11514 9324 11520 9376
rect 11572 9364 11578 9376
rect 12158 9364 12164 9376
rect 11572 9336 12164 9364
rect 11572 9324 11578 9336
rect 12158 9324 12164 9336
rect 12216 9364 12222 9376
rect 18414 9364 18420 9376
rect 12216 9336 18420 9364
rect 12216 9324 12222 9336
rect 18414 9324 18420 9336
rect 18472 9324 18478 9376
rect 22281 9367 22339 9373
rect 22281 9333 22293 9367
rect 22327 9364 22339 9367
rect 22830 9364 22836 9376
rect 22327 9336 22836 9364
rect 22327 9333 22339 9336
rect 22281 9327 22339 9333
rect 22830 9324 22836 9336
rect 22888 9324 22894 9376
rect 1104 9274 25852 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 12214 9274
rect 12266 9222 12278 9274
rect 12330 9222 12342 9274
rect 12394 9222 12406 9274
rect 12458 9222 12470 9274
rect 12522 9222 20214 9274
rect 20266 9222 20278 9274
rect 20330 9222 20342 9274
rect 20394 9222 20406 9274
rect 20458 9222 20470 9274
rect 20522 9222 25852 9274
rect 1104 9200 25852 9222
rect 6546 9120 6552 9172
rect 6604 9120 6610 9172
rect 6730 9120 6736 9172
rect 6788 9160 6794 9172
rect 7101 9163 7159 9169
rect 7101 9160 7113 9163
rect 6788 9132 7113 9160
rect 6788 9120 6794 9132
rect 7101 9129 7113 9132
rect 7147 9129 7159 9163
rect 7101 9123 7159 9129
rect 7929 9163 7987 9169
rect 7929 9129 7941 9163
rect 7975 9160 7987 9163
rect 11057 9163 11115 9169
rect 7975 9132 10640 9160
rect 7975 9129 7987 9132
rect 7929 9123 7987 9129
rect 3513 9095 3571 9101
rect 3513 9061 3525 9095
rect 3559 9092 3571 9095
rect 3970 9092 3976 9104
rect 3559 9064 3976 9092
rect 3559 9061 3571 9064
rect 3513 9055 3571 9061
rect 3970 9052 3976 9064
rect 4028 9092 4034 9104
rect 4065 9095 4123 9101
rect 4065 9092 4077 9095
rect 4028 9064 4077 9092
rect 4028 9052 4034 9064
rect 4065 9061 4077 9064
rect 4111 9061 4123 9095
rect 6089 9095 6147 9101
rect 4065 9055 4123 9061
rect 4264 9064 5948 9092
rect 3145 9027 3203 9033
rect 3145 8993 3157 9027
rect 3191 9024 3203 9027
rect 3234 9024 3240 9036
rect 3191 8996 3240 9024
rect 3191 8993 3203 8996
rect 3145 8987 3203 8993
rect 3234 8984 3240 8996
rect 3292 9024 3298 9036
rect 4264 9024 4292 9064
rect 3292 8996 4292 9024
rect 3292 8984 3298 8996
rect 4614 8984 4620 9036
rect 4672 8984 4678 9036
rect 2222 8916 2228 8968
rect 2280 8916 2286 8968
rect 3329 8959 3387 8965
rect 3329 8925 3341 8959
rect 3375 8956 3387 8959
rect 3602 8956 3608 8968
rect 3375 8928 3608 8956
rect 3375 8925 3387 8928
rect 3329 8919 3387 8925
rect 3602 8916 3608 8928
rect 3660 8916 3666 8968
rect 4706 8916 4712 8968
rect 4764 8916 4770 8968
rect 4982 8916 4988 8968
rect 5040 8956 5046 8968
rect 5736 8965 5764 9064
rect 5813 9027 5871 9033
rect 5813 8993 5825 9027
rect 5859 8993 5871 9027
rect 5920 9024 5948 9064
rect 6089 9061 6101 9095
rect 6135 9092 6147 9095
rect 10612 9092 10640 9132
rect 11057 9129 11069 9163
rect 11103 9160 11115 9163
rect 11146 9160 11152 9172
rect 11103 9132 11152 9160
rect 11103 9129 11115 9132
rect 11057 9123 11115 9129
rect 11146 9120 11152 9132
rect 11204 9120 11210 9172
rect 11256 9132 15332 9160
rect 11256 9092 11284 9132
rect 6135 9064 7052 9092
rect 10612 9064 11284 9092
rect 15197 9095 15255 9101
rect 6135 9061 6147 9064
rect 6089 9055 6147 9061
rect 5920 8996 6500 9024
rect 5813 8987 5871 8993
rect 5077 8959 5135 8965
rect 5077 8956 5089 8959
rect 5040 8928 5089 8956
rect 5040 8916 5046 8928
rect 5077 8925 5089 8928
rect 5123 8925 5135 8959
rect 5077 8919 5135 8925
rect 5721 8959 5779 8965
rect 5721 8925 5733 8959
rect 5767 8925 5779 8959
rect 5828 8956 5856 8987
rect 6472 8965 6500 8996
rect 7024 8965 7052 9064
rect 15197 9061 15209 9095
rect 15243 9061 15255 9095
rect 15304 9092 15332 9132
rect 15470 9120 15476 9172
rect 15528 9120 15534 9172
rect 17678 9120 17684 9172
rect 17736 9120 17742 9172
rect 22094 9120 22100 9172
rect 22152 9160 22158 9172
rect 23385 9163 23443 9169
rect 23385 9160 23397 9163
rect 22152 9132 23397 9160
rect 22152 9120 22158 9132
rect 23385 9129 23397 9132
rect 23431 9129 23443 9163
rect 23385 9123 23443 9129
rect 24394 9120 24400 9172
rect 24452 9160 24458 9172
rect 24489 9163 24547 9169
rect 24489 9160 24501 9163
rect 24452 9132 24501 9160
rect 24452 9120 24458 9132
rect 24489 9129 24501 9132
rect 24535 9129 24547 9163
rect 24489 9123 24547 9129
rect 15304 9064 16436 9092
rect 15197 9055 15255 9061
rect 7834 8984 7840 9036
rect 7892 9024 7898 9036
rect 9309 9027 9367 9033
rect 9309 9024 9321 9027
rect 7892 8996 9321 9024
rect 7892 8984 7898 8996
rect 9309 8993 9321 8996
rect 9355 8993 9367 9027
rect 9309 8987 9367 8993
rect 9582 8984 9588 9036
rect 9640 8984 9646 9036
rect 13170 8984 13176 9036
rect 13228 9024 13234 9036
rect 13449 9027 13507 9033
rect 13449 9024 13461 9027
rect 13228 8996 13461 9024
rect 13228 8984 13234 8996
rect 13449 8993 13461 8996
rect 13495 8993 13507 9027
rect 13449 8987 13507 8993
rect 14550 8984 14556 9036
rect 14608 8984 14614 9036
rect 15212 9024 15240 9055
rect 15212 8996 16160 9024
rect 6365 8959 6423 8965
rect 6365 8956 6377 8959
rect 5828 8928 6377 8956
rect 5721 8919 5779 8925
rect 6365 8925 6377 8928
rect 6411 8925 6423 8959
rect 6365 8919 6423 8925
rect 6458 8959 6516 8965
rect 6458 8925 6470 8959
rect 6504 8925 6516 8959
rect 6458 8919 6516 8925
rect 7009 8959 7067 8965
rect 7009 8925 7021 8959
rect 7055 8925 7067 8959
rect 7009 8919 7067 8925
rect 4065 8891 4123 8897
rect 4065 8857 4077 8891
rect 4111 8888 4123 8891
rect 4724 8888 4752 8916
rect 4111 8860 4752 8888
rect 6380 8888 6408 8919
rect 7098 8916 7104 8968
rect 7156 8956 7162 8968
rect 7193 8959 7251 8965
rect 7193 8956 7205 8959
rect 7156 8928 7205 8956
rect 7156 8916 7162 8928
rect 7193 8925 7205 8928
rect 7239 8925 7251 8959
rect 7193 8919 7251 8925
rect 8018 8916 8024 8968
rect 8076 8956 8082 8968
rect 8113 8959 8171 8965
rect 8113 8956 8125 8959
rect 8076 8928 8125 8956
rect 8076 8916 8082 8928
rect 8113 8925 8125 8928
rect 8159 8925 8171 8959
rect 8113 8919 8171 8925
rect 14737 8959 14795 8965
rect 14737 8925 14749 8959
rect 14783 8956 14795 8959
rect 15286 8956 15292 8968
rect 14783 8928 15292 8956
rect 14783 8925 14795 8928
rect 14737 8919 14795 8925
rect 15286 8916 15292 8928
rect 15344 8916 15350 8968
rect 15378 8916 15384 8968
rect 15436 8956 15442 8968
rect 15473 8959 15531 8965
rect 15473 8956 15485 8959
rect 15436 8928 15485 8956
rect 15436 8916 15442 8928
rect 15473 8925 15485 8928
rect 15519 8925 15531 8959
rect 15473 8919 15531 8925
rect 6380 8860 8064 8888
rect 4111 8857 4123 8860
rect 4065 8851 4123 8857
rect 1762 8780 1768 8832
rect 1820 8820 1826 8832
rect 2041 8823 2099 8829
rect 2041 8820 2053 8823
rect 1820 8792 2053 8820
rect 1820 8780 1826 8792
rect 2041 8789 2053 8792
rect 2087 8789 2099 8823
rect 2041 8783 2099 8789
rect 4522 8780 4528 8832
rect 4580 8780 4586 8832
rect 4706 8780 4712 8832
rect 4764 8820 4770 8832
rect 4801 8823 4859 8829
rect 4801 8820 4813 8823
rect 4764 8792 4813 8820
rect 4764 8780 4770 8792
rect 4801 8789 4813 8792
rect 4847 8789 4859 8823
rect 4801 8783 4859 8789
rect 4890 8780 4896 8832
rect 4948 8820 4954 8832
rect 5169 8823 5227 8829
rect 5169 8820 5181 8823
rect 4948 8792 5181 8820
rect 4948 8780 4954 8792
rect 5169 8789 5181 8792
rect 5215 8789 5227 8823
rect 5169 8783 5227 8789
rect 5994 8780 6000 8832
rect 6052 8820 6058 8832
rect 6089 8823 6147 8829
rect 6089 8820 6101 8823
rect 6052 8792 6101 8820
rect 6052 8780 6058 8792
rect 6089 8789 6101 8792
rect 6135 8789 6147 8823
rect 6089 8783 6147 8789
rect 7282 8780 7288 8832
rect 7340 8820 7346 8832
rect 7929 8823 7987 8829
rect 7929 8820 7941 8823
rect 7340 8792 7941 8820
rect 7340 8780 7346 8792
rect 7929 8789 7941 8792
rect 7975 8789 7987 8823
rect 8036 8820 8064 8860
rect 10594 8848 10600 8900
rect 10652 8848 10658 8900
rect 10888 8860 11744 8888
rect 10888 8820 10916 8860
rect 11716 8832 11744 8860
rect 11882 8848 11888 8900
rect 11940 8888 11946 8900
rect 13173 8891 13231 8897
rect 11940 8860 12006 8888
rect 11940 8848 11946 8860
rect 13173 8857 13185 8891
rect 13219 8857 13231 8891
rect 15488 8888 15516 8919
rect 15654 8916 15660 8968
rect 15712 8916 15718 8968
rect 16132 8965 16160 8996
rect 16117 8959 16175 8965
rect 16117 8925 16129 8959
rect 16163 8925 16175 8959
rect 16117 8919 16175 8925
rect 16022 8888 16028 8900
rect 15488 8860 16028 8888
rect 13173 8851 13231 8857
rect 8036 8792 10916 8820
rect 7929 8783 7987 8789
rect 11698 8780 11704 8832
rect 11756 8780 11762 8832
rect 12434 8780 12440 8832
rect 12492 8820 12498 8832
rect 13188 8820 13216 8851
rect 16022 8848 16028 8860
rect 16080 8888 16086 8900
rect 16408 8888 16436 9064
rect 17218 9052 17224 9104
rect 17276 9092 17282 9104
rect 21361 9095 21419 9101
rect 21361 9092 21373 9095
rect 17276 9064 21373 9092
rect 17276 9052 17282 9064
rect 21361 9061 21373 9064
rect 21407 9061 21419 9095
rect 21361 9055 21419 9061
rect 18414 8984 18420 9036
rect 18472 9024 18478 9036
rect 19797 9027 19855 9033
rect 19797 9024 19809 9027
rect 18472 8996 19809 9024
rect 18472 8984 18478 8996
rect 19797 8993 19809 8996
rect 19843 8993 19855 9027
rect 19797 8987 19855 8993
rect 19978 8984 19984 9036
rect 20036 8984 20042 9036
rect 22830 8984 22836 9036
rect 22888 8984 22894 9036
rect 23106 8984 23112 9036
rect 23164 8984 23170 9036
rect 23382 8984 23388 9036
rect 23440 9024 23446 9036
rect 23937 9027 23995 9033
rect 23937 9024 23949 9027
rect 23440 8996 23949 9024
rect 23440 8984 23446 8996
rect 23937 8993 23949 8996
rect 23983 8993 23995 9027
rect 23937 8987 23995 8993
rect 16482 8916 16488 8968
rect 16540 8958 16546 8968
rect 17681 8959 17739 8965
rect 16540 8956 16574 8958
rect 17681 8956 17693 8959
rect 16540 8928 17693 8956
rect 16540 8916 16546 8928
rect 17681 8925 17693 8928
rect 17727 8925 17739 8959
rect 17681 8919 17739 8925
rect 17865 8959 17923 8965
rect 17865 8925 17877 8959
rect 17911 8956 17923 8959
rect 17954 8956 17960 8968
rect 17911 8928 17960 8956
rect 17911 8925 17923 8928
rect 17865 8919 17923 8925
rect 17494 8888 17500 8900
rect 16080 8860 16252 8888
rect 16408 8860 17500 8888
rect 16080 8848 16086 8860
rect 12492 8792 13216 8820
rect 12492 8780 12498 8792
rect 14826 8780 14832 8832
rect 14884 8780 14890 8832
rect 15470 8780 15476 8832
rect 15528 8820 15534 8832
rect 15933 8823 15991 8829
rect 15933 8820 15945 8823
rect 15528 8792 15945 8820
rect 15528 8780 15534 8792
rect 15933 8789 15945 8792
rect 15979 8789 15991 8823
rect 16224 8820 16252 8860
rect 17494 8848 17500 8860
rect 17552 8848 17558 8900
rect 17696 8888 17724 8919
rect 17954 8916 17960 8928
rect 18012 8916 18018 8968
rect 19705 8959 19763 8965
rect 19705 8925 19717 8959
rect 19751 8956 19763 8959
rect 21450 8956 21456 8968
rect 19751 8928 21456 8956
rect 19751 8925 19763 8928
rect 19705 8919 19763 8925
rect 21450 8916 21456 8928
rect 21508 8916 21514 8968
rect 24118 8916 24124 8968
rect 24176 8956 24182 8968
rect 24489 8959 24547 8965
rect 24489 8956 24501 8959
rect 24176 8928 24501 8956
rect 24176 8916 24182 8928
rect 24489 8925 24501 8928
rect 24535 8925 24547 8959
rect 24489 8919 24547 8925
rect 24673 8959 24731 8965
rect 24673 8925 24685 8959
rect 24719 8925 24731 8959
rect 24673 8919 24731 8925
rect 19150 8888 19156 8900
rect 17696 8860 19156 8888
rect 19150 8848 19156 8860
rect 19208 8848 19214 8900
rect 20070 8848 20076 8900
rect 20128 8888 20134 8900
rect 20533 8891 20591 8897
rect 20533 8888 20545 8891
rect 20128 8860 20545 8888
rect 20128 8848 20134 8860
rect 20533 8857 20545 8860
rect 20579 8857 20591 8891
rect 20533 8851 20591 8857
rect 21818 8848 21824 8900
rect 21876 8848 21882 8900
rect 23474 8848 23480 8900
rect 23532 8888 23538 8900
rect 24688 8888 24716 8919
rect 23532 8860 24716 8888
rect 23532 8848 23538 8860
rect 16482 8820 16488 8832
rect 16224 8792 16488 8820
rect 15933 8783 15991 8789
rect 16482 8780 16488 8792
rect 16540 8780 16546 8832
rect 19337 8823 19395 8829
rect 19337 8789 19349 8823
rect 19383 8820 19395 8823
rect 19518 8820 19524 8832
rect 19383 8792 19524 8820
rect 19383 8789 19395 8792
rect 19337 8783 19395 8789
rect 19518 8780 19524 8792
rect 19576 8780 19582 8832
rect 20622 8780 20628 8832
rect 20680 8780 20686 8832
rect 21361 8823 21419 8829
rect 21361 8789 21373 8823
rect 21407 8820 21419 8823
rect 23753 8823 23811 8829
rect 23753 8820 23765 8823
rect 21407 8792 23765 8820
rect 21407 8789 21419 8792
rect 21361 8783 21419 8789
rect 23753 8789 23765 8792
rect 23799 8789 23811 8823
rect 23753 8783 23811 8789
rect 23845 8823 23903 8829
rect 23845 8789 23857 8823
rect 23891 8820 23903 8823
rect 24118 8820 24124 8832
rect 23891 8792 24124 8820
rect 23891 8789 23903 8792
rect 23845 8783 23903 8789
rect 24118 8780 24124 8792
rect 24176 8780 24182 8832
rect 1104 8730 25852 8752
rect 1104 8678 8214 8730
rect 8266 8678 8278 8730
rect 8330 8678 8342 8730
rect 8394 8678 8406 8730
rect 8458 8678 8470 8730
rect 8522 8678 16214 8730
rect 16266 8678 16278 8730
rect 16330 8678 16342 8730
rect 16394 8678 16406 8730
rect 16458 8678 16470 8730
rect 16522 8678 24214 8730
rect 24266 8678 24278 8730
rect 24330 8678 24342 8730
rect 24394 8678 24406 8730
rect 24458 8678 24470 8730
rect 24522 8678 25852 8730
rect 1104 8656 25852 8678
rect 1302 8576 1308 8628
rect 1360 8616 1366 8628
rect 1360 8588 3556 8616
rect 1360 8576 1366 8588
rect 1762 8508 1768 8560
rect 1820 8508 1826 8560
rect 2774 8508 2780 8560
rect 2832 8508 2838 8560
rect 3528 8489 3556 8588
rect 3602 8576 3608 8628
rect 3660 8576 3666 8628
rect 3878 8576 3884 8628
rect 3936 8616 3942 8628
rect 4065 8619 4123 8625
rect 4065 8616 4077 8619
rect 3936 8588 4077 8616
rect 3936 8576 3942 8588
rect 4065 8585 4077 8588
rect 4111 8585 4123 8619
rect 4065 8579 4123 8585
rect 7098 8576 7104 8628
rect 7156 8616 7162 8628
rect 8294 8616 8300 8628
rect 7156 8588 8300 8616
rect 7156 8576 7162 8588
rect 8294 8576 8300 8588
rect 8352 8616 8358 8628
rect 10045 8619 10103 8625
rect 10045 8616 10057 8619
rect 8352 8588 10057 8616
rect 8352 8576 8358 8588
rect 10045 8585 10057 8588
rect 10091 8585 10103 8619
rect 10045 8579 10103 8585
rect 10410 8576 10416 8628
rect 10468 8576 10474 8628
rect 10594 8576 10600 8628
rect 10652 8616 10658 8628
rect 10781 8619 10839 8625
rect 10781 8616 10793 8619
rect 10652 8588 10793 8616
rect 10652 8576 10658 8588
rect 10781 8585 10793 8588
rect 10827 8585 10839 8619
rect 10781 8579 10839 8585
rect 11882 8576 11888 8628
rect 11940 8576 11946 8628
rect 12434 8576 12440 8628
rect 12492 8576 12498 8628
rect 12713 8619 12771 8625
rect 12713 8585 12725 8619
rect 12759 8585 12771 8619
rect 12713 8579 12771 8585
rect 13173 8619 13231 8625
rect 13173 8585 13185 8619
rect 13219 8616 13231 8619
rect 17218 8616 17224 8628
rect 13219 8588 17224 8616
rect 13219 8585 13231 8588
rect 13173 8579 13231 8585
rect 4617 8551 4675 8557
rect 4617 8517 4629 8551
rect 4663 8548 4675 8551
rect 5074 8548 5080 8560
rect 4663 8520 5080 8548
rect 4663 8517 4675 8520
rect 4617 8511 4675 8517
rect 5074 8508 5080 8520
rect 5132 8508 5138 8560
rect 7374 8508 7380 8560
rect 7432 8548 7438 8560
rect 7469 8551 7527 8557
rect 7469 8548 7481 8551
rect 7432 8520 7481 8548
rect 7432 8508 7438 8520
rect 7469 8517 7481 8520
rect 7515 8517 7527 8551
rect 9309 8551 9367 8557
rect 9309 8548 9321 8551
rect 8694 8520 9321 8548
rect 7469 8511 7527 8517
rect 9309 8517 9321 8520
rect 9355 8517 9367 8551
rect 9309 8511 9367 8517
rect 9953 8551 10011 8557
rect 9953 8517 9965 8551
rect 9999 8548 10011 8551
rect 11514 8548 11520 8560
rect 9999 8520 11520 8548
rect 9999 8517 10011 8520
rect 9953 8511 10011 8517
rect 11514 8508 11520 8520
rect 11572 8508 11578 8560
rect 3513 8483 3571 8489
rect 3513 8449 3525 8483
rect 3559 8449 3571 8483
rect 3513 8443 3571 8449
rect 4062 8440 4068 8492
rect 4120 8480 4126 8492
rect 4341 8483 4399 8489
rect 4341 8480 4353 8483
rect 4120 8452 4353 8480
rect 4120 8440 4126 8452
rect 4341 8449 4353 8452
rect 4387 8449 4399 8483
rect 4798 8480 4804 8492
rect 4341 8443 4399 8449
rect 4632 8452 4804 8480
rect 1486 8372 1492 8424
rect 1544 8372 1550 8424
rect 3234 8372 3240 8424
rect 3292 8372 3298 8424
rect 4229 8415 4287 8421
rect 4229 8381 4241 8415
rect 4275 8412 4287 8415
rect 4632 8412 4660 8452
rect 4798 8440 4804 8452
rect 4856 8480 4862 8492
rect 4985 8483 5043 8489
rect 4985 8480 4997 8483
rect 4856 8452 4997 8480
rect 4856 8440 4862 8452
rect 4985 8449 4997 8452
rect 5031 8449 5043 8483
rect 4985 8443 5043 8449
rect 5166 8440 5172 8492
rect 5224 8440 5230 8492
rect 5261 8483 5319 8489
rect 5261 8449 5273 8483
rect 5307 8449 5319 8483
rect 5261 8443 5319 8449
rect 5905 8483 5963 8489
rect 5905 8449 5917 8483
rect 5951 8480 5963 8483
rect 7098 8480 7104 8492
rect 5951 8452 7104 8480
rect 5951 8449 5963 8452
rect 5905 8443 5963 8449
rect 4275 8384 4660 8412
rect 4275 8381 4287 8384
rect 4229 8375 4287 8381
rect 4706 8372 4712 8424
rect 4764 8372 4770 8424
rect 4890 8372 4896 8424
rect 4948 8412 4954 8424
rect 5276 8412 5304 8443
rect 7098 8440 7104 8452
rect 7156 8440 7162 8492
rect 7190 8440 7196 8492
rect 7248 8440 7254 8492
rect 9217 8483 9275 8489
rect 9217 8449 9229 8483
rect 9263 8449 9275 8483
rect 9217 8443 9275 8449
rect 9401 8483 9459 8489
rect 9401 8449 9413 8483
rect 9447 8480 9459 8483
rect 9674 8480 9680 8492
rect 9447 8452 9680 8480
rect 9447 8449 9459 8452
rect 9401 8443 9459 8449
rect 4948 8384 5304 8412
rect 4948 8372 4954 8384
rect 5994 8372 6000 8424
rect 6052 8372 6058 8424
rect 9232 8412 9260 8443
rect 9674 8440 9680 8452
rect 9732 8480 9738 8492
rect 10689 8483 10747 8489
rect 9732 8452 10640 8480
rect 9732 8440 9738 8452
rect 10612 8424 10640 8452
rect 10689 8449 10701 8483
rect 10735 8480 10747 8483
rect 10778 8480 10784 8492
rect 10735 8452 10784 8480
rect 10735 8449 10747 8452
rect 10689 8443 10747 8449
rect 10778 8440 10784 8452
rect 10836 8440 10842 8492
rect 10873 8483 10931 8489
rect 10873 8449 10885 8483
rect 10919 8449 10931 8483
rect 10873 8443 10931 8449
rect 9306 8412 9312 8424
rect 9232 8384 9312 8412
rect 9306 8372 9312 8384
rect 9364 8372 9370 8424
rect 9766 8372 9772 8424
rect 9824 8372 9830 8424
rect 10594 8372 10600 8424
rect 10652 8412 10658 8424
rect 10888 8412 10916 8443
rect 11238 8440 11244 8492
rect 11296 8480 11302 8492
rect 11793 8483 11851 8489
rect 11793 8480 11805 8483
rect 11296 8452 11805 8480
rect 11296 8440 11302 8452
rect 11793 8449 11805 8452
rect 11839 8480 11851 8483
rect 11882 8480 11888 8492
rect 11839 8452 11888 8480
rect 11839 8449 11851 8452
rect 11793 8443 11851 8449
rect 11882 8440 11888 8452
rect 11940 8440 11946 8492
rect 11974 8440 11980 8492
rect 12032 8440 12038 8492
rect 12253 8483 12311 8489
rect 12253 8449 12265 8483
rect 12299 8480 12311 8483
rect 12728 8480 12756 8579
rect 17218 8576 17224 8588
rect 17276 8576 17282 8628
rect 17313 8619 17371 8625
rect 17313 8585 17325 8619
rect 17359 8585 17371 8619
rect 17313 8579 17371 8585
rect 15010 8508 15016 8560
rect 15068 8508 15074 8560
rect 15470 8508 15476 8560
rect 15528 8508 15534 8560
rect 12299 8452 12756 8480
rect 13081 8483 13139 8489
rect 12299 8449 12311 8452
rect 12253 8443 12311 8449
rect 13081 8449 13093 8483
rect 13127 8449 13139 8483
rect 13081 8443 13139 8449
rect 17037 8483 17095 8489
rect 17037 8449 17049 8483
rect 17083 8480 17095 8483
rect 17328 8480 17356 8579
rect 17770 8576 17776 8628
rect 17828 8576 17834 8628
rect 18690 8576 18696 8628
rect 18748 8576 18754 8628
rect 19705 8619 19763 8625
rect 19705 8585 19717 8619
rect 19751 8616 19763 8619
rect 19794 8616 19800 8628
rect 19751 8588 19800 8616
rect 19751 8585 19763 8588
rect 19705 8579 19763 8585
rect 19794 8576 19800 8588
rect 19852 8576 19858 8628
rect 20441 8619 20499 8625
rect 20441 8585 20453 8619
rect 20487 8616 20499 8619
rect 20898 8616 20904 8628
rect 20487 8588 20904 8616
rect 20487 8585 20499 8588
rect 20441 8579 20499 8585
rect 20898 8576 20904 8588
rect 20956 8576 20962 8628
rect 21818 8576 21824 8628
rect 21876 8616 21882 8628
rect 22005 8619 22063 8625
rect 22005 8616 22017 8619
rect 21876 8588 22017 8616
rect 21876 8576 21882 8588
rect 22005 8585 22017 8588
rect 22051 8585 22063 8619
rect 22005 8579 22063 8585
rect 18966 8508 18972 8560
rect 19024 8548 19030 8560
rect 19242 8548 19248 8560
rect 19024 8520 19248 8548
rect 19024 8508 19030 8520
rect 19242 8508 19248 8520
rect 19300 8548 19306 8560
rect 20622 8548 20628 8560
rect 19300 8520 20628 8548
rect 19300 8508 19306 8520
rect 17083 8452 17356 8480
rect 17083 8449 17095 8452
rect 17037 8443 17095 8449
rect 10652 8384 10916 8412
rect 10652 8372 10658 8384
rect 11698 8372 11704 8424
rect 11756 8412 11762 8424
rect 13096 8412 13124 8443
rect 17586 8440 17592 8492
rect 17644 8480 17650 8492
rect 17681 8483 17739 8489
rect 17681 8480 17693 8483
rect 17644 8452 17693 8480
rect 17644 8440 17650 8452
rect 17681 8449 17693 8452
rect 17727 8449 17739 8483
rect 17681 8443 17739 8449
rect 18782 8440 18788 8492
rect 18840 8440 18846 8492
rect 19518 8440 19524 8492
rect 19576 8440 19582 8492
rect 20364 8489 20392 8520
rect 20622 8508 20628 8520
rect 20680 8548 20686 8560
rect 20680 8520 21496 8548
rect 20680 8508 20686 8520
rect 20349 8483 20407 8489
rect 20349 8449 20361 8483
rect 20395 8449 20407 8483
rect 20349 8443 20407 8449
rect 20533 8483 20591 8489
rect 20533 8449 20545 8483
rect 20579 8449 20591 8483
rect 20533 8443 20591 8449
rect 11756 8384 13124 8412
rect 13357 8415 13415 8421
rect 11756 8372 11762 8384
rect 13357 8381 13369 8415
rect 13403 8381 13415 8415
rect 13357 8375 13415 8381
rect 14001 8415 14059 8421
rect 14001 8381 14013 8415
rect 14047 8412 14059 8415
rect 14826 8412 14832 8424
rect 14047 8384 14832 8412
rect 14047 8381 14059 8384
rect 14001 8375 14059 8381
rect 4522 8304 4528 8356
rect 4580 8344 4586 8356
rect 4985 8347 5043 8353
rect 4985 8344 4997 8347
rect 4580 8316 4997 8344
rect 4580 8304 4586 8316
rect 4985 8313 4997 8316
rect 5031 8313 5043 8347
rect 4985 8307 5043 8313
rect 5534 8304 5540 8356
rect 5592 8304 5598 8356
rect 8754 8304 8760 8356
rect 8812 8344 8818 8356
rect 8941 8347 8999 8353
rect 8941 8344 8953 8347
rect 8812 8316 8953 8344
rect 8812 8304 8818 8316
rect 8941 8313 8953 8316
rect 8987 8313 8999 8347
rect 13372 8344 13400 8375
rect 14826 8372 14832 8384
rect 14884 8372 14890 8424
rect 15749 8415 15807 8421
rect 15749 8381 15761 8415
rect 15795 8412 15807 8415
rect 16666 8412 16672 8424
rect 15795 8384 16672 8412
rect 15795 8381 15807 8384
rect 15749 8375 15807 8381
rect 16666 8372 16672 8384
rect 16724 8372 16730 8424
rect 17494 8372 17500 8424
rect 17552 8412 17558 8424
rect 17957 8415 18015 8421
rect 17957 8412 17969 8415
rect 17552 8384 17969 8412
rect 17552 8372 17558 8384
rect 17957 8381 17969 8384
rect 18003 8412 18015 8415
rect 18601 8415 18659 8421
rect 18601 8412 18613 8415
rect 18003 8384 18613 8412
rect 18003 8381 18015 8384
rect 17957 8375 18015 8381
rect 18601 8381 18613 8384
rect 18647 8412 18659 8415
rect 18647 8384 19564 8412
rect 18647 8381 18659 8384
rect 18601 8375 18659 8381
rect 13814 8344 13820 8356
rect 13372 8316 13820 8344
rect 8941 8307 8999 8313
rect 13814 8304 13820 8316
rect 13872 8344 13878 8356
rect 14458 8344 14464 8356
rect 13872 8316 14464 8344
rect 13872 8304 13878 8316
rect 14458 8304 14464 8316
rect 14516 8304 14522 8356
rect 19153 8347 19211 8353
rect 19153 8313 19165 8347
rect 19199 8344 19211 8347
rect 19426 8344 19432 8356
rect 19199 8316 19432 8344
rect 19199 8313 19211 8316
rect 19153 8307 19211 8313
rect 19426 8304 19432 8316
rect 19484 8304 19490 8356
rect 19536 8344 19564 8384
rect 19610 8372 19616 8424
rect 19668 8412 19674 8424
rect 20548 8412 20576 8443
rect 20806 8440 20812 8492
rect 20864 8440 20870 8492
rect 21468 8489 21496 8520
rect 23566 8508 23572 8560
rect 23624 8548 23630 8560
rect 23624 8520 24150 8548
rect 23624 8508 23630 8520
rect 21269 8483 21327 8489
rect 21269 8449 21281 8483
rect 21315 8449 21327 8483
rect 21269 8443 21327 8449
rect 21453 8483 21511 8489
rect 21453 8449 21465 8483
rect 21499 8449 21511 8483
rect 21453 8443 21511 8449
rect 21284 8412 21312 8443
rect 19668 8384 21312 8412
rect 21468 8412 21496 8443
rect 21818 8440 21824 8492
rect 21876 8480 21882 8492
rect 21913 8483 21971 8489
rect 21913 8480 21925 8483
rect 21876 8452 21925 8480
rect 21876 8440 21882 8452
rect 21913 8449 21925 8452
rect 21959 8449 21971 8483
rect 21913 8443 21971 8449
rect 22097 8483 22155 8489
rect 22097 8449 22109 8483
rect 22143 8449 22155 8483
rect 22097 8443 22155 8449
rect 22002 8412 22008 8424
rect 21468 8384 22008 8412
rect 19668 8372 19674 8384
rect 22002 8372 22008 8384
rect 22060 8372 22066 8424
rect 19536 8316 20024 8344
rect 16853 8279 16911 8285
rect 16853 8245 16865 8279
rect 16899 8276 16911 8279
rect 16942 8276 16948 8288
rect 16899 8248 16948 8276
rect 16899 8245 16911 8248
rect 16853 8239 16911 8245
rect 16942 8236 16948 8248
rect 17000 8236 17006 8288
rect 19996 8276 20024 8316
rect 20070 8304 20076 8356
rect 20128 8344 20134 8356
rect 22112 8344 22140 8443
rect 23106 8440 23112 8492
rect 23164 8480 23170 8492
rect 23385 8483 23443 8489
rect 23385 8480 23397 8483
rect 23164 8452 23397 8480
rect 23164 8440 23170 8452
rect 23385 8449 23397 8452
rect 23431 8449 23443 8483
rect 23385 8443 23443 8449
rect 23658 8372 23664 8424
rect 23716 8372 23722 8424
rect 20128 8316 23520 8344
rect 20128 8304 20134 8316
rect 23492 8288 23520 8316
rect 20714 8276 20720 8288
rect 19996 8248 20720 8276
rect 20714 8236 20720 8248
rect 20772 8236 20778 8288
rect 20990 8236 20996 8288
rect 21048 8236 21054 8288
rect 21269 8279 21327 8285
rect 21269 8245 21281 8279
rect 21315 8276 21327 8279
rect 22922 8276 22928 8288
rect 21315 8248 22928 8276
rect 21315 8245 21327 8248
rect 21269 8239 21327 8245
rect 22922 8236 22928 8248
rect 22980 8236 22986 8288
rect 23474 8236 23480 8288
rect 23532 8236 23538 8288
rect 25130 8236 25136 8288
rect 25188 8236 25194 8288
rect 1104 8186 25852 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 12214 8186
rect 12266 8134 12278 8186
rect 12330 8134 12342 8186
rect 12394 8134 12406 8186
rect 12458 8134 12470 8186
rect 12522 8134 20214 8186
rect 20266 8134 20278 8186
rect 20330 8134 20342 8186
rect 20394 8134 20406 8186
rect 20458 8134 20470 8186
rect 20522 8134 25852 8186
rect 1104 8112 25852 8134
rect 2222 8032 2228 8084
rect 2280 8072 2286 8084
rect 2593 8075 2651 8081
rect 2593 8072 2605 8075
rect 2280 8044 2605 8072
rect 2280 8032 2286 8044
rect 2593 8041 2605 8044
rect 2639 8041 2651 8075
rect 2593 8035 2651 8041
rect 3602 8032 3608 8084
rect 3660 8072 3666 8084
rect 4065 8075 4123 8081
rect 4065 8072 4077 8075
rect 3660 8044 4077 8072
rect 3660 8032 3666 8044
rect 4065 8041 4077 8044
rect 4111 8041 4123 8075
rect 4065 8035 4123 8041
rect 4525 8075 4583 8081
rect 4525 8041 4537 8075
rect 4571 8072 4583 8075
rect 4614 8072 4620 8084
rect 4571 8044 4620 8072
rect 4571 8041 4583 8044
rect 4525 8035 4583 8041
rect 4614 8032 4620 8044
rect 4672 8032 4678 8084
rect 6089 8075 6147 8081
rect 5092 8044 6040 8072
rect 2317 8007 2375 8013
rect 2317 7973 2329 8007
rect 2363 8004 2375 8007
rect 2774 8004 2780 8016
rect 2363 7976 2780 8004
rect 2363 7973 2375 7976
rect 2317 7967 2375 7973
rect 2774 7964 2780 7976
rect 2832 7964 2838 8016
rect 5092 8004 5120 8044
rect 3068 7976 5120 8004
rect 2498 7936 2504 7948
rect 2148 7908 2504 7936
rect 2148 7877 2176 7908
rect 2498 7896 2504 7908
rect 2556 7936 2562 7948
rect 3068 7936 3096 7976
rect 5166 7964 5172 8016
rect 5224 7964 5230 8016
rect 5537 8007 5595 8013
rect 5537 7973 5549 8007
rect 5583 7973 5595 8007
rect 6012 8004 6040 8044
rect 6089 8041 6101 8075
rect 6135 8072 6147 8075
rect 6362 8072 6368 8084
rect 6135 8044 6368 8072
rect 6135 8041 6147 8044
rect 6089 8035 6147 8041
rect 6362 8032 6368 8044
rect 6420 8032 6426 8084
rect 10686 8032 10692 8084
rect 10744 8032 10750 8084
rect 11882 8032 11888 8084
rect 11940 8072 11946 8084
rect 12250 8072 12256 8084
rect 11940 8044 12256 8072
rect 11940 8032 11946 8044
rect 12250 8032 12256 8044
rect 12308 8072 12314 8084
rect 12437 8075 12495 8081
rect 12437 8072 12449 8075
rect 12308 8044 12449 8072
rect 12308 8032 12314 8044
rect 12437 8041 12449 8044
rect 12483 8041 12495 8075
rect 12437 8035 12495 8041
rect 14369 8075 14427 8081
rect 14369 8041 14381 8075
rect 14415 8072 14427 8075
rect 14550 8072 14556 8084
rect 14415 8044 14556 8072
rect 14415 8041 14427 8044
rect 14369 8035 14427 8041
rect 14550 8032 14556 8044
rect 14608 8032 14614 8084
rect 15010 8032 15016 8084
rect 15068 8072 15074 8084
rect 15381 8075 15439 8081
rect 15381 8072 15393 8075
rect 15068 8044 15393 8072
rect 15068 8032 15074 8044
rect 15381 8041 15393 8044
rect 15427 8041 15439 8075
rect 18230 8072 18236 8084
rect 15381 8035 15439 8041
rect 16546 8044 18236 8072
rect 9674 8004 9680 8016
rect 6012 7976 9680 8004
rect 5537 7967 5595 7973
rect 2556 7908 3096 7936
rect 3145 7939 3203 7945
rect 2556 7896 2562 7908
rect 3145 7905 3157 7939
rect 3191 7936 3203 7939
rect 3418 7936 3424 7948
rect 3191 7908 3424 7936
rect 3191 7905 3203 7908
rect 3145 7899 3203 7905
rect 3418 7896 3424 7908
rect 3476 7896 3482 7948
rect 5184 7936 5212 7964
rect 4264 7908 5212 7936
rect 5552 7936 5580 7967
rect 9674 7964 9680 7976
rect 9732 7964 9738 8016
rect 12360 7976 15516 8004
rect 8205 7939 8263 7945
rect 8205 7936 8217 7939
rect 5552 7908 6132 7936
rect 2133 7871 2191 7877
rect 2133 7837 2145 7871
rect 2179 7837 2191 7871
rect 2133 7831 2191 7837
rect 2317 7871 2375 7877
rect 2317 7837 2329 7871
rect 2363 7868 2375 7871
rect 2682 7868 2688 7880
rect 2363 7840 2688 7868
rect 2363 7837 2375 7840
rect 2317 7831 2375 7837
rect 2682 7828 2688 7840
rect 2740 7828 2746 7880
rect 2961 7871 3019 7877
rect 2961 7837 2973 7871
rect 3007 7868 3019 7871
rect 3234 7868 3240 7880
rect 3007 7840 3240 7868
rect 3007 7837 3019 7840
rect 2961 7831 3019 7837
rect 3234 7828 3240 7840
rect 3292 7868 3298 7880
rect 3973 7871 4031 7877
rect 3973 7868 3985 7871
rect 3292 7840 3985 7868
rect 3292 7828 3298 7840
rect 3973 7837 3985 7840
rect 4019 7837 4031 7871
rect 3973 7831 4031 7837
rect 4062 7828 4068 7880
rect 4120 7868 4126 7880
rect 4264 7877 4292 7908
rect 4249 7871 4307 7877
rect 4249 7868 4261 7871
rect 4120 7840 4261 7868
rect 4120 7828 4126 7840
rect 4249 7837 4261 7840
rect 4295 7837 4307 7871
rect 4249 7831 4307 7837
rect 4341 7871 4399 7877
rect 4341 7837 4353 7871
rect 4387 7868 4399 7871
rect 4890 7868 4896 7880
rect 4387 7840 4896 7868
rect 4387 7837 4399 7840
rect 4341 7831 4399 7837
rect 4890 7828 4896 7840
rect 4948 7828 4954 7880
rect 5168 7871 5226 7877
rect 5168 7837 5180 7871
rect 5214 7837 5226 7871
rect 5168 7831 5226 7837
rect 5261 7871 5319 7877
rect 5261 7837 5273 7871
rect 5307 7868 5319 7871
rect 5552 7868 5580 7908
rect 5307 7840 5580 7868
rect 5307 7837 5319 7840
rect 5261 7831 5319 7837
rect 3053 7735 3111 7741
rect 3053 7701 3065 7735
rect 3099 7732 3111 7735
rect 4430 7732 4436 7744
rect 3099 7704 4436 7732
rect 3099 7701 3111 7704
rect 3053 7695 3111 7701
rect 4430 7692 4436 7704
rect 4488 7692 4494 7744
rect 4890 7692 4896 7744
rect 4948 7692 4954 7744
rect 5184 7732 5212 7831
rect 5810 7828 5816 7880
rect 5868 7828 5874 7880
rect 6104 7877 6132 7908
rect 7944 7908 8217 7936
rect 6089 7871 6147 7877
rect 6089 7837 6101 7871
rect 6135 7837 6147 7871
rect 6089 7831 6147 7837
rect 6362 7828 6368 7880
rect 6420 7828 6426 7880
rect 7444 7871 7502 7877
rect 7444 7837 7456 7871
rect 7490 7868 7502 7871
rect 7944 7868 7972 7908
rect 8205 7905 8217 7908
rect 8251 7936 8263 7939
rect 8570 7936 8576 7948
rect 8251 7908 8576 7936
rect 8251 7905 8263 7908
rect 8205 7899 8263 7905
rect 8570 7896 8576 7908
rect 8628 7896 8634 7948
rect 9766 7896 9772 7948
rect 9824 7936 9830 7948
rect 10045 7939 10103 7945
rect 10045 7936 10057 7939
rect 9824 7908 10057 7936
rect 9824 7896 9830 7908
rect 10045 7905 10057 7908
rect 10091 7905 10103 7939
rect 10045 7899 10103 7905
rect 10229 7939 10287 7945
rect 10229 7905 10241 7939
rect 10275 7936 10287 7939
rect 11146 7936 11152 7948
rect 10275 7908 11152 7936
rect 10275 7905 10287 7908
rect 10229 7899 10287 7905
rect 11146 7896 11152 7908
rect 11204 7896 11210 7948
rect 7490 7840 7972 7868
rect 8021 7871 8079 7877
rect 7490 7837 7502 7840
rect 7444 7831 7502 7837
rect 8021 7837 8033 7871
rect 8067 7868 8079 7871
rect 8110 7868 8116 7880
rect 8067 7840 8116 7868
rect 8067 7837 8079 7840
rect 8021 7831 8079 7837
rect 8110 7828 8116 7840
rect 8168 7828 8174 7880
rect 8294 7828 8300 7880
rect 8352 7868 8358 7880
rect 8662 7868 8668 7880
rect 8352 7840 8668 7868
rect 8352 7828 8358 7840
rect 8662 7828 8668 7840
rect 8720 7828 8726 7880
rect 12066 7828 12072 7880
rect 12124 7868 12130 7880
rect 12360 7877 12388 7976
rect 12309 7871 12388 7877
rect 12309 7868 12321 7871
rect 12124 7840 12321 7868
rect 12124 7828 12130 7840
rect 12309 7837 12321 7840
rect 12355 7840 12388 7871
rect 12529 7871 12587 7877
rect 12355 7837 12367 7840
rect 12309 7831 12367 7837
rect 12529 7837 12541 7871
rect 12575 7868 12587 7871
rect 12805 7871 12863 7877
rect 12805 7868 12817 7871
rect 12575 7840 12817 7868
rect 12575 7837 12587 7840
rect 12529 7831 12587 7837
rect 12805 7837 12817 7840
rect 12851 7837 12863 7871
rect 12805 7831 12863 7837
rect 12989 7871 13047 7877
rect 12989 7837 13001 7871
rect 13035 7837 13047 7871
rect 12989 7831 13047 7837
rect 5534 7760 5540 7812
rect 5592 7760 5598 7812
rect 5994 7800 6000 7812
rect 5644 7772 6000 7800
rect 5644 7732 5672 7772
rect 5994 7760 6000 7772
rect 6052 7800 6058 7812
rect 6273 7803 6331 7809
rect 6273 7800 6285 7803
rect 6052 7772 6285 7800
rect 6052 7760 6058 7772
rect 6273 7769 6285 7772
rect 6319 7769 6331 7803
rect 6273 7763 6331 7769
rect 9493 7803 9551 7809
rect 9493 7769 9505 7803
rect 9539 7800 9551 7803
rect 10134 7800 10140 7812
rect 9539 7772 10140 7800
rect 9539 7769 9551 7772
rect 9493 7763 9551 7769
rect 10134 7760 10140 7772
rect 10192 7760 10198 7812
rect 11790 7760 11796 7812
rect 11848 7800 11854 7812
rect 13004 7800 13032 7831
rect 14182 7828 14188 7880
rect 14240 7828 14246 7880
rect 14734 7828 14740 7880
rect 14792 7868 14798 7880
rect 14921 7871 14979 7877
rect 14921 7868 14933 7871
rect 14792 7840 14933 7868
rect 14792 7828 14798 7840
rect 14921 7837 14933 7840
rect 14967 7837 14979 7871
rect 14921 7831 14979 7837
rect 15381 7871 15439 7877
rect 15381 7837 15393 7871
rect 15427 7837 15439 7871
rect 15488 7868 15516 7976
rect 15565 7871 15623 7877
rect 15565 7868 15577 7871
rect 15488 7840 15577 7868
rect 15381 7831 15439 7837
rect 15565 7837 15577 7840
rect 15611 7868 15623 7871
rect 15654 7868 15660 7880
rect 15611 7840 15660 7868
rect 15611 7837 15623 7840
rect 15565 7831 15623 7837
rect 11848 7772 13032 7800
rect 15105 7803 15163 7809
rect 11848 7760 11854 7772
rect 15105 7769 15117 7803
rect 15151 7800 15163 7803
rect 15194 7800 15200 7812
rect 15151 7772 15200 7800
rect 15151 7769 15163 7772
rect 15105 7763 15163 7769
rect 15194 7760 15200 7772
rect 15252 7760 15258 7812
rect 15396 7800 15424 7831
rect 15654 7828 15660 7840
rect 15712 7868 15718 7880
rect 15841 7871 15899 7877
rect 15841 7868 15853 7871
rect 15712 7840 15853 7868
rect 15712 7828 15718 7840
rect 15841 7837 15853 7840
rect 15887 7837 15899 7871
rect 15841 7831 15899 7837
rect 16022 7828 16028 7880
rect 16080 7828 16086 7880
rect 16546 7800 16574 8044
rect 18230 8032 18236 8044
rect 18288 8072 18294 8084
rect 23385 8075 23443 8081
rect 18288 8044 18736 8072
rect 18288 8032 18294 8044
rect 16942 7896 16948 7948
rect 17000 7896 17006 7948
rect 16666 7828 16672 7880
rect 16724 7828 16730 7880
rect 18708 7877 18736 8044
rect 23385 8041 23397 8075
rect 23431 8072 23443 8075
rect 23566 8072 23572 8084
rect 23431 8044 23572 8072
rect 23431 8041 23443 8044
rect 23385 8035 23443 8041
rect 23566 8032 23572 8044
rect 23624 8032 23630 8084
rect 23658 8032 23664 8084
rect 23716 8072 23722 8084
rect 23845 8075 23903 8081
rect 23845 8072 23857 8075
rect 23716 8044 23857 8072
rect 23716 8032 23722 8044
rect 23845 8041 23857 8044
rect 23891 8041 23903 8075
rect 23845 8035 23903 8041
rect 24026 8032 24032 8084
rect 24084 8072 24090 8084
rect 24084 8044 24992 8072
rect 24084 8032 24090 8044
rect 23106 7964 23112 8016
rect 23164 7964 23170 8016
rect 24489 8007 24547 8013
rect 24489 7973 24501 8007
rect 24535 7973 24547 8007
rect 24964 8004 24992 8044
rect 24964 7976 25084 8004
rect 24489 7967 24547 7973
rect 20990 7896 20996 7948
rect 21048 7936 21054 7948
rect 21453 7939 21511 7945
rect 21453 7936 21465 7939
rect 21048 7908 21465 7936
rect 21048 7896 21054 7908
rect 21453 7905 21465 7908
rect 21499 7905 21511 7939
rect 21453 7899 21511 7905
rect 21729 7939 21787 7945
rect 21729 7905 21741 7939
rect 21775 7936 21787 7939
rect 22370 7936 22376 7948
rect 21775 7908 22376 7936
rect 21775 7905 21787 7908
rect 21729 7899 21787 7905
rect 22370 7896 22376 7908
rect 22428 7936 22434 7948
rect 23124 7936 23152 7964
rect 22428 7908 23152 7936
rect 22428 7896 22434 7908
rect 18693 7871 18751 7877
rect 18693 7837 18705 7871
rect 18739 7837 18751 7871
rect 18693 7831 18751 7837
rect 18877 7871 18935 7877
rect 18877 7837 18889 7871
rect 18923 7868 18935 7871
rect 18966 7868 18972 7880
rect 18923 7840 18972 7868
rect 18923 7837 18935 7840
rect 18877 7831 18935 7837
rect 18966 7828 18972 7840
rect 19024 7828 19030 7880
rect 19426 7828 19432 7880
rect 19484 7868 19490 7880
rect 19521 7871 19579 7877
rect 19521 7868 19533 7871
rect 19484 7840 19533 7868
rect 19484 7828 19490 7840
rect 19521 7837 19533 7840
rect 19567 7837 19579 7871
rect 19521 7831 19579 7837
rect 20346 7828 20352 7880
rect 20404 7828 20410 7880
rect 23106 7828 23112 7880
rect 23164 7828 23170 7880
rect 23385 7871 23443 7877
rect 23385 7837 23397 7871
rect 23431 7837 23443 7871
rect 23385 7831 23443 7837
rect 18785 7803 18843 7809
rect 18785 7800 18797 7803
rect 15396 7772 16574 7800
rect 18170 7772 18797 7800
rect 5184 7704 5672 7732
rect 5718 7692 5724 7744
rect 5776 7692 5782 7744
rect 7515 7735 7573 7741
rect 7515 7701 7527 7735
rect 7561 7732 7573 7735
rect 7742 7732 7748 7744
rect 7561 7704 7748 7732
rect 7561 7701 7573 7704
rect 7515 7695 7573 7701
rect 7742 7692 7748 7704
rect 7800 7692 7806 7744
rect 7837 7735 7895 7741
rect 7837 7701 7849 7735
rect 7883 7732 7895 7735
rect 8018 7732 8024 7744
rect 7883 7704 8024 7732
rect 7883 7701 7895 7704
rect 7837 7695 7895 7701
rect 8018 7692 8024 7704
rect 8076 7692 8082 7744
rect 8938 7692 8944 7744
rect 8996 7732 9002 7744
rect 10321 7735 10379 7741
rect 10321 7732 10333 7735
rect 8996 7704 10333 7732
rect 8996 7692 9002 7704
rect 10321 7701 10333 7704
rect 10367 7701 10379 7735
rect 10321 7695 10379 7701
rect 12894 7692 12900 7744
rect 12952 7692 12958 7744
rect 13630 7692 13636 7744
rect 13688 7732 13694 7744
rect 15396 7732 15424 7772
rect 18785 7769 18797 7772
rect 18831 7769 18843 7803
rect 18785 7763 18843 7769
rect 22554 7760 22560 7812
rect 22612 7800 22618 7812
rect 23400 7800 23428 7831
rect 23474 7828 23480 7880
rect 23532 7868 23538 7880
rect 23569 7871 23627 7877
rect 23569 7868 23581 7871
rect 23532 7840 23581 7868
rect 23532 7828 23538 7840
rect 23569 7837 23581 7840
rect 23615 7837 23627 7871
rect 23569 7831 23627 7837
rect 24029 7871 24087 7877
rect 24029 7837 24041 7871
rect 24075 7868 24087 7871
rect 24504 7868 24532 7967
rect 24762 7896 24768 7948
rect 24820 7936 24826 7948
rect 25056 7945 25084 7976
rect 24949 7939 25007 7945
rect 24949 7936 24961 7939
rect 24820 7908 24961 7936
rect 24820 7896 24826 7908
rect 24949 7905 24961 7908
rect 24995 7905 25007 7939
rect 24949 7899 25007 7905
rect 25041 7939 25099 7945
rect 25041 7905 25053 7939
rect 25087 7905 25099 7939
rect 25041 7899 25099 7905
rect 24075 7840 24532 7868
rect 24857 7871 24915 7877
rect 24075 7837 24087 7840
rect 24029 7831 24087 7837
rect 24857 7837 24869 7871
rect 24903 7868 24915 7871
rect 25130 7868 25136 7880
rect 24903 7840 25136 7868
rect 24903 7837 24915 7840
rect 24857 7831 24915 7837
rect 25130 7828 25136 7840
rect 25188 7828 25194 7880
rect 22612 7772 23428 7800
rect 22612 7760 22618 7772
rect 13688 7704 15424 7732
rect 13688 7692 13694 7704
rect 15838 7692 15844 7744
rect 15896 7732 15902 7744
rect 15933 7735 15991 7741
rect 15933 7732 15945 7735
rect 15896 7704 15945 7732
rect 15896 7692 15902 7704
rect 15933 7701 15945 7704
rect 15979 7701 15991 7735
rect 15933 7695 15991 7701
rect 17586 7692 17592 7744
rect 17644 7732 17650 7744
rect 18417 7735 18475 7741
rect 18417 7732 18429 7735
rect 17644 7704 18429 7732
rect 17644 7692 17650 7704
rect 18417 7701 18429 7704
rect 18463 7701 18475 7735
rect 18417 7695 18475 7701
rect 18874 7692 18880 7744
rect 18932 7732 18938 7744
rect 19337 7735 19395 7741
rect 19337 7732 19349 7735
rect 18932 7704 19349 7732
rect 18932 7692 18938 7704
rect 19337 7701 19349 7704
rect 19383 7701 19395 7735
rect 19337 7695 19395 7701
rect 19981 7735 20039 7741
rect 19981 7701 19993 7735
rect 20027 7732 20039 7735
rect 21082 7732 21088 7744
rect 20027 7704 21088 7732
rect 20027 7701 20039 7704
rect 19981 7695 20039 7701
rect 21082 7692 21088 7704
rect 21140 7692 21146 7744
rect 22646 7692 22652 7744
rect 22704 7732 22710 7744
rect 22925 7735 22983 7741
rect 22925 7732 22937 7735
rect 22704 7704 22937 7732
rect 22704 7692 22710 7704
rect 22925 7701 22937 7704
rect 22971 7701 22983 7735
rect 22925 7695 22983 7701
rect 1104 7642 25852 7664
rect 1104 7590 8214 7642
rect 8266 7590 8278 7642
rect 8330 7590 8342 7642
rect 8394 7590 8406 7642
rect 8458 7590 8470 7642
rect 8522 7590 16214 7642
rect 16266 7590 16278 7642
rect 16330 7590 16342 7642
rect 16394 7590 16406 7642
rect 16458 7590 16470 7642
rect 16522 7590 24214 7642
rect 24266 7590 24278 7642
rect 24330 7590 24342 7642
rect 24394 7590 24406 7642
rect 24458 7590 24470 7642
rect 24522 7590 25852 7642
rect 1104 7568 25852 7590
rect 4430 7488 4436 7540
rect 4488 7488 4494 7540
rect 5718 7528 5724 7540
rect 4724 7500 5724 7528
rect 3789 7463 3847 7469
rect 3789 7429 3801 7463
rect 3835 7460 3847 7463
rect 4724 7460 4752 7500
rect 5718 7488 5724 7500
rect 5776 7488 5782 7540
rect 5810 7488 5816 7540
rect 5868 7528 5874 7540
rect 6086 7528 6092 7540
rect 5868 7500 6092 7528
rect 5868 7488 5874 7500
rect 6086 7488 6092 7500
rect 6144 7528 6150 7540
rect 6549 7531 6607 7537
rect 6549 7528 6561 7531
rect 6144 7500 6561 7528
rect 6144 7488 6150 7500
rect 6549 7497 6561 7500
rect 6595 7497 6607 7531
rect 6549 7491 6607 7497
rect 7098 7488 7104 7540
rect 7156 7488 7162 7540
rect 11054 7528 11060 7540
rect 7208 7500 11060 7528
rect 4890 7460 4896 7472
rect 3835 7432 4752 7460
rect 4815 7432 4896 7460
rect 3835 7429 3847 7432
rect 3789 7423 3847 7429
rect 1854 7352 1860 7404
rect 1912 7392 1918 7404
rect 2498 7392 2504 7404
rect 1912 7364 2504 7392
rect 1912 7352 1918 7364
rect 2498 7352 2504 7364
rect 2556 7352 2562 7404
rect 2682 7352 2688 7404
rect 2740 7352 2746 7404
rect 4062 7392 4068 7404
rect 4023 7364 4068 7392
rect 4062 7352 4068 7364
rect 4120 7352 4126 7404
rect 4815 7401 4843 7432
rect 4890 7420 4896 7432
rect 4948 7420 4954 7472
rect 6270 7460 6276 7472
rect 5092 7432 6276 7460
rect 4157 7395 4215 7401
rect 4157 7361 4169 7395
rect 4203 7361 4215 7395
rect 4157 7355 4215 7361
rect 4775 7395 4843 7401
rect 4775 7361 4787 7395
rect 4821 7364 4843 7395
rect 4821 7361 4833 7364
rect 4775 7355 4833 7361
rect 4172 7256 4200 7355
rect 4893 7327 4951 7333
rect 4893 7293 4905 7327
rect 4939 7324 4951 7327
rect 5092 7324 5120 7432
rect 6270 7420 6276 7432
rect 6328 7420 6334 7472
rect 7208 7460 7236 7500
rect 11054 7488 11060 7500
rect 11112 7488 11118 7540
rect 13630 7528 13636 7540
rect 12084 7500 13636 7528
rect 6380 7432 7236 7460
rect 5166 7352 5172 7404
rect 5224 7392 5230 7404
rect 5445 7395 5503 7401
rect 5445 7392 5457 7395
rect 5224 7364 5457 7392
rect 5224 7352 5230 7364
rect 5445 7361 5457 7364
rect 5491 7361 5503 7395
rect 5445 7355 5503 7361
rect 4939 7296 5120 7324
rect 5353 7327 5411 7333
rect 4939 7293 4951 7296
rect 4893 7287 4951 7293
rect 5353 7293 5365 7327
rect 5399 7324 5411 7327
rect 6380 7324 6408 7432
rect 8018 7420 8024 7472
rect 8076 7420 8082 7472
rect 9582 7460 9588 7472
rect 9246 7432 9588 7460
rect 9582 7420 9588 7432
rect 9640 7420 9646 7472
rect 6457 7395 6515 7401
rect 6457 7361 6469 7395
rect 6503 7361 6515 7395
rect 6457 7355 6515 7361
rect 5399 7296 6408 7324
rect 5399 7293 5411 7296
rect 5353 7287 5411 7293
rect 5368 7256 5396 7287
rect 4172 7228 5396 7256
rect 5534 7216 5540 7268
rect 5592 7256 5598 7268
rect 5813 7259 5871 7265
rect 5813 7256 5825 7259
rect 5592 7228 5825 7256
rect 5592 7216 5598 7228
rect 5813 7225 5825 7228
rect 5859 7256 5871 7259
rect 6472 7256 6500 7355
rect 6638 7352 6644 7404
rect 6696 7352 6702 7404
rect 7006 7352 7012 7404
rect 7064 7352 7070 7404
rect 7285 7395 7343 7401
rect 7285 7392 7297 7395
rect 7116 7364 7297 7392
rect 6656 7324 6684 7352
rect 7116 7324 7144 7364
rect 7285 7361 7297 7364
rect 7331 7361 7343 7395
rect 7285 7355 7343 7361
rect 9769 7395 9827 7401
rect 9769 7361 9781 7395
rect 9815 7392 9827 7395
rect 10134 7392 10140 7404
rect 9815 7364 10140 7392
rect 9815 7361 9827 7364
rect 9769 7355 9827 7361
rect 10134 7352 10140 7364
rect 10192 7352 10198 7404
rect 11790 7352 11796 7404
rect 11848 7352 11854 7404
rect 11974 7352 11980 7404
rect 12032 7392 12038 7404
rect 12084 7401 12112 7500
rect 13630 7488 13636 7500
rect 13688 7488 13694 7540
rect 14182 7488 14188 7540
rect 14240 7528 14246 7540
rect 14240 7500 14780 7528
rect 14240 7488 14246 7500
rect 12894 7420 12900 7472
rect 12952 7460 12958 7472
rect 14752 7460 14780 7500
rect 16666 7488 16672 7540
rect 16724 7528 16730 7540
rect 16724 7500 19196 7528
rect 16724 7488 16730 7500
rect 15102 7460 15108 7472
rect 12952 7432 13938 7460
rect 14752 7432 15108 7460
rect 12952 7420 12958 7432
rect 15102 7420 15108 7432
rect 15160 7460 15166 7472
rect 16761 7463 16819 7469
rect 16761 7460 16773 7463
rect 15160 7432 16773 7460
rect 15160 7420 15166 7432
rect 16761 7429 16773 7432
rect 16807 7429 16819 7463
rect 16761 7423 16819 7429
rect 18874 7420 18880 7472
rect 18932 7420 18938 7472
rect 12069 7395 12127 7401
rect 12069 7392 12081 7395
rect 12032 7364 12081 7392
rect 12032 7352 12038 7364
rect 12069 7361 12081 7364
rect 12115 7361 12127 7395
rect 12069 7355 12127 7361
rect 12250 7352 12256 7404
rect 12308 7352 12314 7404
rect 15473 7395 15531 7401
rect 15473 7361 15485 7395
rect 15519 7392 15531 7395
rect 15654 7392 15660 7404
rect 15519 7364 15660 7392
rect 15519 7361 15531 7364
rect 15473 7355 15531 7361
rect 15654 7352 15660 7364
rect 15712 7352 15718 7404
rect 16942 7352 16948 7404
rect 17000 7352 17006 7404
rect 17770 7352 17776 7404
rect 17828 7352 17834 7404
rect 19168 7401 19196 7500
rect 20346 7488 20352 7540
rect 20404 7488 20410 7540
rect 20717 7531 20775 7537
rect 20717 7497 20729 7531
rect 20763 7528 20775 7531
rect 20806 7528 20812 7540
rect 20763 7500 20812 7528
rect 20763 7497 20775 7500
rect 20717 7491 20775 7497
rect 20806 7488 20812 7500
rect 20864 7488 20870 7540
rect 21082 7488 21088 7540
rect 21140 7488 21146 7540
rect 21177 7531 21235 7537
rect 21177 7497 21189 7531
rect 21223 7528 21235 7531
rect 21910 7528 21916 7540
rect 21223 7500 21916 7528
rect 21223 7497 21235 7500
rect 21177 7491 21235 7497
rect 21910 7488 21916 7500
rect 21968 7488 21974 7540
rect 24118 7488 24124 7540
rect 24176 7488 24182 7540
rect 19426 7420 19432 7472
rect 19484 7460 19490 7472
rect 22554 7460 22560 7472
rect 19484 7432 22560 7460
rect 19484 7420 19490 7432
rect 19153 7395 19211 7401
rect 19153 7361 19165 7395
rect 19199 7361 19211 7395
rect 19153 7355 19211 7361
rect 19242 7352 19248 7404
rect 19300 7392 19306 7404
rect 19705 7395 19763 7401
rect 19705 7392 19717 7395
rect 19300 7364 19717 7392
rect 19300 7352 19306 7364
rect 19705 7361 19717 7364
rect 19751 7361 19763 7395
rect 19705 7355 19763 7361
rect 19889 7395 19947 7401
rect 19889 7361 19901 7395
rect 19935 7392 19947 7395
rect 20070 7392 20076 7404
rect 19935 7364 20076 7392
rect 19935 7361 19947 7364
rect 19889 7355 19947 7361
rect 20070 7352 20076 7364
rect 20128 7392 20134 7404
rect 20456 7401 20484 7432
rect 22554 7420 22560 7432
rect 22612 7420 22618 7472
rect 22646 7420 22652 7472
rect 22704 7420 22710 7472
rect 22922 7420 22928 7472
rect 22980 7460 22986 7472
rect 22980 7432 23138 7460
rect 22980 7420 22986 7432
rect 20257 7395 20315 7401
rect 20257 7392 20269 7395
rect 20128 7364 20269 7392
rect 20128 7352 20134 7364
rect 20257 7361 20269 7364
rect 20303 7361 20315 7395
rect 20257 7355 20315 7361
rect 20441 7395 20499 7401
rect 20441 7361 20453 7395
rect 20487 7361 20499 7395
rect 20441 7355 20499 7361
rect 21818 7352 21824 7404
rect 21876 7392 21882 7404
rect 21913 7395 21971 7401
rect 21913 7392 21925 7395
rect 21876 7364 21925 7392
rect 21876 7352 21882 7364
rect 21913 7361 21925 7364
rect 21959 7361 21971 7395
rect 21913 7355 21971 7361
rect 22002 7352 22008 7404
rect 22060 7392 22066 7404
rect 22097 7395 22155 7401
rect 22097 7392 22109 7395
rect 22060 7364 22109 7392
rect 22060 7352 22066 7364
rect 22097 7361 22109 7364
rect 22143 7361 22155 7395
rect 22097 7355 22155 7361
rect 22370 7352 22376 7404
rect 22428 7352 22434 7404
rect 24578 7352 24584 7404
rect 24636 7352 24642 7404
rect 6656 7296 7144 7324
rect 7190 7284 7196 7336
rect 7248 7324 7254 7336
rect 7745 7327 7803 7333
rect 7745 7324 7757 7327
rect 7248 7296 7757 7324
rect 7248 7284 7254 7296
rect 7745 7293 7757 7296
rect 7791 7324 7803 7327
rect 9030 7324 9036 7336
rect 7791 7296 9036 7324
rect 7791 7293 7803 7296
rect 7745 7287 7803 7293
rect 9030 7284 9036 7296
rect 9088 7284 9094 7336
rect 13170 7284 13176 7336
rect 13228 7284 13234 7336
rect 13446 7284 13452 7336
rect 13504 7284 13510 7336
rect 15197 7327 15255 7333
rect 15197 7293 15209 7327
rect 15243 7324 15255 7327
rect 15378 7324 15384 7336
rect 15243 7296 15384 7324
rect 15243 7293 15255 7296
rect 15197 7287 15255 7293
rect 15378 7284 15384 7296
rect 15436 7284 15442 7336
rect 17405 7327 17463 7333
rect 17405 7293 17417 7327
rect 17451 7324 17463 7327
rect 18782 7324 18788 7336
rect 17451 7296 18788 7324
rect 17451 7293 17463 7296
rect 17405 7287 17463 7293
rect 18782 7284 18788 7296
rect 18840 7284 18846 7336
rect 20714 7284 20720 7336
rect 20772 7324 20778 7336
rect 21361 7327 21419 7333
rect 21361 7324 21373 7327
rect 20772 7296 21373 7324
rect 20772 7284 20778 7296
rect 21361 7293 21373 7296
rect 21407 7324 21419 7327
rect 24026 7324 24032 7336
rect 21407 7296 24032 7324
rect 21407 7293 21419 7296
rect 21361 7287 21419 7293
rect 24026 7284 24032 7296
rect 24084 7284 24090 7336
rect 5859 7228 6500 7256
rect 5859 7225 5871 7228
rect 5813 7219 5871 7225
rect 23934 7216 23940 7268
rect 23992 7256 23998 7268
rect 24397 7259 24455 7265
rect 24397 7256 24409 7259
rect 23992 7228 24409 7256
rect 23992 7216 23998 7228
rect 24397 7225 24409 7228
rect 24443 7225 24455 7259
rect 24397 7219 24455 7225
rect 2685 7191 2743 7197
rect 2685 7157 2697 7191
rect 2731 7188 2743 7191
rect 2774 7188 2780 7200
rect 2731 7160 2780 7188
rect 2731 7157 2743 7160
rect 2685 7151 2743 7157
rect 2774 7148 2780 7160
rect 2832 7148 2838 7200
rect 7466 7148 7472 7200
rect 7524 7148 7530 7200
rect 9490 7148 9496 7200
rect 9548 7148 9554 7200
rect 9950 7148 9956 7200
rect 10008 7148 10014 7200
rect 11606 7148 11612 7200
rect 11664 7148 11670 7200
rect 11974 7148 11980 7200
rect 12032 7188 12038 7200
rect 12069 7191 12127 7197
rect 12069 7188 12081 7191
rect 12032 7160 12081 7188
rect 12032 7148 12038 7160
rect 12069 7157 12081 7160
rect 12115 7157 12127 7191
rect 12069 7151 12127 7157
rect 14918 7148 14924 7200
rect 14976 7148 14982 7200
rect 21910 7148 21916 7200
rect 21968 7148 21974 7200
rect 1104 7098 25852 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 12214 7098
rect 12266 7046 12278 7098
rect 12330 7046 12342 7098
rect 12394 7046 12406 7098
rect 12458 7046 12470 7098
rect 12522 7046 20214 7098
rect 20266 7046 20278 7098
rect 20330 7046 20342 7098
rect 20394 7046 20406 7098
rect 20458 7046 20470 7098
rect 20522 7046 25852 7098
rect 1104 7024 25852 7046
rect 3237 6987 3295 6993
rect 3237 6953 3249 6987
rect 3283 6984 3295 6987
rect 4062 6984 4068 6996
rect 3283 6956 4068 6984
rect 3283 6953 3295 6956
rect 3237 6947 3295 6953
rect 4062 6944 4068 6956
rect 4120 6944 4126 6996
rect 5994 6944 6000 6996
rect 6052 6944 6058 6996
rect 7098 6944 7104 6996
rect 7156 6984 7162 6996
rect 8481 6987 8539 6993
rect 8481 6984 8493 6987
rect 7156 6956 8493 6984
rect 7156 6944 7162 6956
rect 8481 6953 8493 6956
rect 8527 6984 8539 6987
rect 9217 6987 9275 6993
rect 8527 6956 8892 6984
rect 8527 6953 8539 6956
rect 8481 6947 8539 6953
rect 6638 6916 6644 6928
rect 5368 6888 6644 6916
rect 1486 6808 1492 6860
rect 1544 6808 1550 6860
rect 5166 6848 5172 6860
rect 4448 6820 5172 6848
rect 4448 6789 4476 6820
rect 5166 6808 5172 6820
rect 5224 6808 5230 6860
rect 5368 6789 5396 6888
rect 6638 6876 6644 6888
rect 6696 6916 6702 6928
rect 8754 6916 8760 6928
rect 6696 6888 8760 6916
rect 6696 6876 6702 6888
rect 8754 6876 8760 6888
rect 8812 6876 8818 6928
rect 8864 6916 8892 6956
rect 9217 6953 9229 6987
rect 9263 6984 9275 6987
rect 9766 6984 9772 6996
rect 9263 6956 9772 6984
rect 9263 6953 9275 6956
rect 9217 6947 9275 6953
rect 9766 6944 9772 6956
rect 9824 6944 9830 6996
rect 11228 6987 11286 6993
rect 11228 6953 11240 6987
rect 11274 6984 11286 6987
rect 11606 6984 11612 6996
rect 11274 6956 11612 6984
rect 11274 6953 11286 6956
rect 11228 6947 11286 6953
rect 11606 6944 11612 6956
rect 11664 6944 11670 6996
rect 13446 6944 13452 6996
rect 13504 6984 13510 6996
rect 13633 6987 13691 6993
rect 13633 6984 13645 6987
rect 13504 6956 13645 6984
rect 13504 6944 13510 6956
rect 13633 6953 13645 6956
rect 13679 6953 13691 6987
rect 13633 6947 13691 6953
rect 18509 6987 18567 6993
rect 18509 6953 18521 6987
rect 18555 6984 18567 6987
rect 18598 6984 18604 6996
rect 18555 6956 18604 6984
rect 18555 6953 18567 6956
rect 18509 6947 18567 6953
rect 18598 6944 18604 6956
rect 18656 6984 18662 6996
rect 19242 6984 19248 6996
rect 18656 6956 19248 6984
rect 18656 6944 18662 6956
rect 19242 6944 19248 6956
rect 19300 6944 19306 6996
rect 19518 6944 19524 6996
rect 19576 6984 19582 6996
rect 22370 6984 22376 6996
rect 19576 6956 22376 6984
rect 19576 6944 19582 6956
rect 22370 6944 22376 6956
rect 22428 6944 22434 6996
rect 23106 6944 23112 6996
rect 23164 6984 23170 6996
rect 23201 6987 23259 6993
rect 23201 6984 23213 6987
rect 23164 6956 23213 6984
rect 23164 6944 23170 6956
rect 23201 6953 23213 6956
rect 23247 6953 23259 6987
rect 23201 6947 23259 6953
rect 24489 6987 24547 6993
rect 24489 6953 24501 6987
rect 24535 6984 24547 6987
rect 24578 6984 24584 6996
rect 24535 6956 24584 6984
rect 24535 6953 24547 6956
rect 24489 6947 24547 6953
rect 24578 6944 24584 6956
rect 24636 6944 24642 6996
rect 9398 6916 9404 6928
rect 8864 6888 9404 6916
rect 9398 6876 9404 6888
rect 9456 6876 9462 6928
rect 13170 6916 13176 6928
rect 12360 6888 13176 6916
rect 5445 6851 5503 6857
rect 5445 6817 5457 6851
rect 5491 6848 5503 6851
rect 5534 6848 5540 6860
rect 5491 6820 5540 6848
rect 5491 6817 5503 6820
rect 5445 6811 5503 6817
rect 5534 6808 5540 6820
rect 5592 6808 5598 6860
rect 7374 6808 7380 6860
rect 7432 6808 7438 6860
rect 7466 6808 7472 6860
rect 7524 6848 7530 6860
rect 8662 6848 8668 6860
rect 7524 6820 7880 6848
rect 7524 6808 7530 6820
rect 4433 6783 4491 6789
rect 4433 6749 4445 6783
rect 4479 6749 4491 6783
rect 4433 6743 4491 6749
rect 4709 6783 4767 6789
rect 4709 6749 4721 6783
rect 4755 6780 4767 6783
rect 5353 6783 5411 6789
rect 4755 6752 5120 6780
rect 4755 6749 4767 6752
rect 4709 6743 4767 6749
rect 1762 6672 1768 6724
rect 1820 6672 1826 6724
rect 2774 6672 2780 6724
rect 2832 6672 2838 6724
rect 4617 6715 4675 6721
rect 4617 6681 4629 6715
rect 4663 6712 4675 6715
rect 4798 6712 4804 6724
rect 4663 6684 4804 6712
rect 4663 6681 4675 6684
rect 4617 6675 4675 6681
rect 4798 6672 4804 6684
rect 4856 6672 4862 6724
rect 3142 6604 3148 6656
rect 3200 6644 3206 6656
rect 3237 6647 3295 6653
rect 3237 6644 3249 6647
rect 3200 6616 3249 6644
rect 3200 6604 3206 6616
rect 3237 6613 3249 6616
rect 3283 6613 3295 6647
rect 3237 6607 3295 6613
rect 4709 6647 4767 6653
rect 4709 6613 4721 6647
rect 4755 6644 4767 6647
rect 4890 6644 4896 6656
rect 4755 6616 4896 6644
rect 4755 6613 4767 6616
rect 4709 6607 4767 6613
rect 4890 6604 4896 6616
rect 4948 6604 4954 6656
rect 4985 6647 5043 6653
rect 4985 6613 4997 6647
rect 5031 6644 5043 6647
rect 5092 6644 5120 6752
rect 5353 6749 5365 6783
rect 5399 6749 5411 6783
rect 5353 6743 5411 6749
rect 5626 6740 5632 6792
rect 5684 6780 5690 6792
rect 5813 6783 5871 6789
rect 5813 6780 5825 6783
rect 5684 6752 5825 6780
rect 5684 6740 5690 6752
rect 5813 6749 5825 6752
rect 5859 6749 5871 6783
rect 5813 6743 5871 6749
rect 6086 6740 6092 6792
rect 6144 6740 6150 6792
rect 7653 6783 7711 6789
rect 7653 6749 7665 6783
rect 7699 6749 7711 6783
rect 7653 6743 7711 6749
rect 5718 6672 5724 6724
rect 5776 6712 5782 6724
rect 5905 6715 5963 6721
rect 5905 6712 5917 6715
rect 5776 6684 5917 6712
rect 5776 6672 5782 6684
rect 5905 6681 5917 6684
rect 5951 6681 5963 6715
rect 7668 6712 7696 6743
rect 7742 6740 7748 6792
rect 7800 6740 7806 6792
rect 7852 6789 7880 6820
rect 7944 6820 8668 6848
rect 7837 6783 7895 6789
rect 7837 6749 7849 6783
rect 7883 6749 7895 6783
rect 7837 6743 7895 6749
rect 7944 6712 7972 6820
rect 8662 6808 8668 6820
rect 8720 6848 8726 6860
rect 9490 6848 9496 6860
rect 8720 6820 9496 6848
rect 8720 6808 8726 6820
rect 8018 6740 8024 6792
rect 8076 6740 8082 6792
rect 8570 6780 8576 6792
rect 8312 6752 8576 6780
rect 7668 6684 7972 6712
rect 5905 6675 5963 6681
rect 5442 6644 5448 6656
rect 5031 6616 5448 6644
rect 5031 6613 5043 6616
rect 4985 6607 5043 6613
rect 5442 6604 5448 6616
rect 5500 6604 5506 6656
rect 6086 6604 6092 6656
rect 6144 6644 6150 6656
rect 7098 6644 7104 6656
rect 6144 6616 7104 6644
rect 6144 6604 6150 6616
rect 7098 6604 7104 6616
rect 7156 6604 7162 6656
rect 8312 6653 8340 6752
rect 8570 6740 8576 6752
rect 8628 6780 8634 6792
rect 8628 6752 8800 6780
rect 8628 6740 8634 6752
rect 8662 6672 8668 6724
rect 8720 6672 8726 6724
rect 8772 6712 8800 6752
rect 9416 6721 9444 6820
rect 9490 6808 9496 6820
rect 9548 6808 9554 6860
rect 9582 6808 9588 6860
rect 9640 6848 9646 6860
rect 9769 6851 9827 6857
rect 9769 6848 9781 6851
rect 9640 6820 9781 6848
rect 9640 6808 9646 6820
rect 9769 6817 9781 6820
rect 9815 6817 9827 6851
rect 9769 6811 9827 6817
rect 10962 6808 10968 6860
rect 11020 6848 11026 6860
rect 12360 6848 12388 6888
rect 13170 6876 13176 6888
rect 13228 6876 13234 6928
rect 17954 6876 17960 6928
rect 18012 6916 18018 6928
rect 18966 6916 18972 6928
rect 18012 6888 18972 6916
rect 18012 6876 18018 6888
rect 18966 6876 18972 6888
rect 19024 6876 19030 6928
rect 11020 6820 12388 6848
rect 11020 6808 11026 6820
rect 12434 6808 12440 6860
rect 12492 6848 12498 6860
rect 15013 6851 15071 6857
rect 15013 6848 15025 6851
rect 12492 6820 15025 6848
rect 12492 6808 12498 6820
rect 15013 6817 15025 6820
rect 15059 6848 15071 6851
rect 17126 6848 17132 6860
rect 15059 6820 17132 6848
rect 15059 6817 15071 6820
rect 15013 6811 15071 6817
rect 17126 6808 17132 6820
rect 17184 6808 17190 6860
rect 20625 6851 20683 6857
rect 20625 6817 20637 6851
rect 20671 6848 20683 6851
rect 21358 6848 21364 6860
rect 20671 6820 21364 6848
rect 20671 6817 20683 6820
rect 20625 6811 20683 6817
rect 21358 6808 21364 6820
rect 21416 6808 21422 6860
rect 22646 6808 22652 6860
rect 22704 6848 22710 6860
rect 23753 6851 23811 6857
rect 23753 6848 23765 6851
rect 22704 6820 23765 6848
rect 22704 6808 22710 6820
rect 23753 6817 23765 6820
rect 23799 6817 23811 6851
rect 23753 6811 23811 6817
rect 24946 6808 24952 6860
rect 25004 6848 25010 6860
rect 25041 6851 25099 6857
rect 25041 6848 25053 6851
rect 25004 6820 25053 6848
rect 25004 6808 25010 6820
rect 25041 6817 25053 6820
rect 25087 6817 25099 6851
rect 25041 6811 25099 6817
rect 9677 6783 9735 6789
rect 9677 6780 9689 6783
rect 9600 6752 9689 6780
rect 9185 6715 9243 6721
rect 9185 6712 9197 6715
rect 8772 6684 9197 6712
rect 9185 6681 9197 6684
rect 9231 6681 9243 6715
rect 9185 6675 9243 6681
rect 9401 6715 9459 6721
rect 9401 6681 9413 6715
rect 9447 6681 9459 6715
rect 9401 6675 9459 6681
rect 8297 6647 8355 6653
rect 8297 6613 8309 6647
rect 8343 6613 8355 6647
rect 8297 6607 8355 6613
rect 8465 6647 8523 6653
rect 8465 6613 8477 6647
rect 8511 6644 8523 6647
rect 8570 6644 8576 6656
rect 8511 6616 8576 6644
rect 8511 6613 8523 6616
rect 8465 6607 8523 6613
rect 8570 6604 8576 6616
rect 8628 6604 8634 6656
rect 8846 6604 8852 6656
rect 8904 6644 8910 6656
rect 9033 6647 9091 6653
rect 9033 6644 9045 6647
rect 8904 6616 9045 6644
rect 8904 6604 8910 6616
rect 9033 6613 9045 6616
rect 9079 6613 9091 6647
rect 9033 6607 9091 6613
rect 9306 6604 9312 6656
rect 9364 6644 9370 6656
rect 9600 6644 9628 6752
rect 9677 6749 9689 6752
rect 9723 6749 9735 6783
rect 9677 6743 9735 6749
rect 9861 6783 9919 6789
rect 9861 6749 9873 6783
rect 9907 6780 9919 6783
rect 9950 6780 9956 6792
rect 9907 6752 9956 6780
rect 9907 6749 9919 6752
rect 9861 6743 9919 6749
rect 9950 6740 9956 6752
rect 10008 6740 10014 6792
rect 12618 6740 12624 6792
rect 12676 6780 12682 6792
rect 12989 6783 13047 6789
rect 12989 6780 13001 6783
rect 12676 6752 13001 6780
rect 12676 6740 12682 6752
rect 12989 6749 13001 6752
rect 13035 6749 13047 6783
rect 12989 6743 13047 6749
rect 13817 6783 13875 6789
rect 13817 6749 13829 6783
rect 13863 6749 13875 6783
rect 13817 6743 13875 6749
rect 11974 6672 11980 6724
rect 12032 6672 12038 6724
rect 9364 6616 9628 6644
rect 9364 6604 9370 6616
rect 11054 6604 11060 6656
rect 11112 6644 11118 6656
rect 12250 6644 12256 6656
rect 11112 6616 12256 6644
rect 11112 6604 11118 6616
rect 12250 6604 12256 6616
rect 12308 6644 12314 6656
rect 12713 6647 12771 6653
rect 12713 6644 12725 6647
rect 12308 6616 12725 6644
rect 12308 6604 12314 6616
rect 12713 6613 12725 6616
rect 12759 6613 12771 6647
rect 12713 6607 12771 6613
rect 13173 6647 13231 6653
rect 13173 6613 13185 6647
rect 13219 6644 13231 6647
rect 13722 6644 13728 6656
rect 13219 6616 13728 6644
rect 13219 6613 13231 6616
rect 13173 6607 13231 6613
rect 13722 6604 13728 6616
rect 13780 6604 13786 6656
rect 13832 6644 13860 6743
rect 14826 6740 14832 6792
rect 14884 6740 14890 6792
rect 15654 6740 15660 6792
rect 15712 6780 15718 6792
rect 17865 6783 17923 6789
rect 15712 6752 16574 6780
rect 15712 6740 15718 6752
rect 16546 6712 16574 6752
rect 17865 6749 17877 6783
rect 17911 6780 17923 6783
rect 17954 6780 17960 6792
rect 17911 6752 17960 6780
rect 17911 6749 17923 6752
rect 17865 6743 17923 6749
rect 17954 6740 17960 6752
rect 18012 6740 18018 6792
rect 18049 6783 18107 6789
rect 18049 6749 18061 6783
rect 18095 6780 18107 6783
rect 18230 6780 18236 6792
rect 18095 6752 18236 6780
rect 18095 6749 18107 6752
rect 18049 6743 18107 6749
rect 18230 6740 18236 6752
rect 18288 6740 18294 6792
rect 18325 6783 18383 6789
rect 18325 6749 18337 6783
rect 18371 6749 18383 6783
rect 18325 6743 18383 6749
rect 18340 6712 18368 6743
rect 19518 6740 19524 6792
rect 19576 6780 19582 6792
rect 20349 6783 20407 6789
rect 20349 6780 20361 6783
rect 19576 6752 20361 6780
rect 19576 6740 19582 6752
rect 20349 6749 20361 6752
rect 20395 6749 20407 6783
rect 20349 6743 20407 6749
rect 23569 6783 23627 6789
rect 23569 6749 23581 6783
rect 23615 6780 23627 6783
rect 24118 6780 24124 6792
rect 23615 6752 24124 6780
rect 23615 6749 23627 6752
rect 23569 6743 23627 6749
rect 24118 6740 24124 6752
rect 24176 6740 24182 6792
rect 24857 6783 24915 6789
rect 24857 6749 24869 6783
rect 24903 6780 24915 6783
rect 25130 6780 25136 6792
rect 24903 6752 25136 6780
rect 24903 6749 24915 6752
rect 24857 6743 24915 6749
rect 25130 6740 25136 6752
rect 25188 6740 25194 6792
rect 21910 6712 21916 6724
rect 16546 6684 18368 6712
rect 21850 6684 21916 6712
rect 21910 6672 21916 6684
rect 21968 6672 21974 6724
rect 14461 6647 14519 6653
rect 14461 6644 14473 6647
rect 13832 6616 14473 6644
rect 14461 6613 14473 6616
rect 14507 6613 14519 6647
rect 14461 6607 14519 6613
rect 14918 6604 14924 6656
rect 14976 6604 14982 6656
rect 15470 6604 15476 6656
rect 15528 6604 15534 6656
rect 17770 6604 17776 6656
rect 17828 6644 17834 6656
rect 17957 6647 18015 6653
rect 17957 6644 17969 6647
rect 17828 6616 17969 6644
rect 17828 6604 17834 6616
rect 17957 6613 17969 6616
rect 18003 6613 18015 6647
rect 17957 6607 18015 6613
rect 22094 6604 22100 6656
rect 22152 6604 22158 6656
rect 23661 6647 23719 6653
rect 23661 6613 23673 6647
rect 23707 6644 23719 6647
rect 24949 6647 25007 6653
rect 24949 6644 24961 6647
rect 23707 6616 24961 6644
rect 23707 6613 23719 6616
rect 23661 6607 23719 6613
rect 24949 6613 24961 6616
rect 24995 6644 25007 6647
rect 25038 6644 25044 6656
rect 24995 6616 25044 6644
rect 24995 6613 25007 6616
rect 24949 6607 25007 6613
rect 25038 6604 25044 6616
rect 25096 6604 25102 6656
rect 1104 6554 25852 6576
rect 1104 6502 8214 6554
rect 8266 6502 8278 6554
rect 8330 6502 8342 6554
rect 8394 6502 8406 6554
rect 8458 6502 8470 6554
rect 8522 6502 16214 6554
rect 16266 6502 16278 6554
rect 16330 6502 16342 6554
rect 16394 6502 16406 6554
rect 16458 6502 16470 6554
rect 16522 6502 24214 6554
rect 24266 6502 24278 6554
rect 24330 6502 24342 6554
rect 24394 6502 24406 6554
rect 24458 6502 24470 6554
rect 24522 6502 25852 6554
rect 1104 6480 25852 6502
rect 1762 6400 1768 6452
rect 1820 6440 1826 6452
rect 2133 6443 2191 6449
rect 2133 6440 2145 6443
rect 1820 6412 2145 6440
rect 1820 6400 1826 6412
rect 2133 6409 2145 6412
rect 2179 6409 2191 6443
rect 2133 6403 2191 6409
rect 2777 6443 2835 6449
rect 2777 6409 2789 6443
rect 2823 6409 2835 6443
rect 2777 6403 2835 6409
rect 2317 6307 2375 6313
rect 2317 6273 2329 6307
rect 2363 6304 2375 6307
rect 2792 6304 2820 6403
rect 3142 6400 3148 6452
rect 3200 6400 3206 6452
rect 4724 6412 6224 6440
rect 4724 6313 4752 6412
rect 4798 6332 4804 6384
rect 4856 6332 4862 6384
rect 4890 6332 4896 6384
rect 4948 6372 4954 6384
rect 4948 6344 5948 6372
rect 4948 6332 4954 6344
rect 2363 6276 2820 6304
rect 4709 6307 4767 6313
rect 2363 6273 2375 6276
rect 2317 6267 2375 6273
rect 4709 6273 4721 6307
rect 4755 6273 4767 6307
rect 4816 6304 4844 6332
rect 4816 6276 4936 6304
rect 4709 6267 4767 6273
rect 3237 6239 3295 6245
rect 3237 6205 3249 6239
rect 3283 6205 3295 6239
rect 3237 6199 3295 6205
rect 3252 6168 3280 6199
rect 3418 6196 3424 6248
rect 3476 6236 3482 6248
rect 3970 6236 3976 6248
rect 3476 6208 3976 6236
rect 3476 6196 3482 6208
rect 3970 6196 3976 6208
rect 4028 6196 4034 6248
rect 4801 6239 4859 6245
rect 4801 6205 4813 6239
rect 4847 6205 4859 6239
rect 4908 6236 4936 6276
rect 5166 6264 5172 6316
rect 5224 6264 5230 6316
rect 5261 6307 5319 6313
rect 5261 6273 5273 6307
rect 5307 6273 5319 6307
rect 5261 6267 5319 6273
rect 5276 6236 5304 6267
rect 5442 6264 5448 6316
rect 5500 6264 5506 6316
rect 5920 6313 5948 6344
rect 5905 6307 5963 6313
rect 5905 6273 5917 6307
rect 5951 6273 5963 6307
rect 5905 6267 5963 6273
rect 6089 6307 6147 6313
rect 6089 6273 6101 6307
rect 6135 6273 6147 6307
rect 6196 6304 6224 6412
rect 6362 6400 6368 6452
rect 6420 6440 6426 6452
rect 6457 6443 6515 6449
rect 6457 6440 6469 6443
rect 6420 6412 6469 6440
rect 6420 6400 6426 6412
rect 6457 6409 6469 6412
rect 6503 6409 6515 6443
rect 6457 6403 6515 6409
rect 7006 6400 7012 6452
rect 7064 6440 7070 6452
rect 8113 6443 8171 6449
rect 8113 6440 8125 6443
rect 7064 6412 8125 6440
rect 7064 6400 7070 6412
rect 6733 6307 6791 6313
rect 6733 6304 6745 6307
rect 6196 6276 6745 6304
rect 6089 6267 6147 6273
rect 6733 6273 6745 6276
rect 6779 6304 6791 6307
rect 7098 6304 7104 6316
rect 6779 6276 7104 6304
rect 6779 6273 6791 6276
rect 6733 6267 6791 6273
rect 5534 6236 5540 6248
rect 4908 6208 5540 6236
rect 4801 6199 4859 6205
rect 4341 6171 4399 6177
rect 4341 6168 4353 6171
rect 3252 6140 4353 6168
rect 4341 6137 4353 6140
rect 4387 6137 4399 6171
rect 4816 6168 4844 6199
rect 5534 6196 5540 6208
rect 5592 6196 5598 6248
rect 5629 6239 5687 6245
rect 5629 6205 5641 6239
rect 5675 6236 5687 6239
rect 6104 6236 6132 6267
rect 7098 6264 7104 6276
rect 7156 6264 7162 6316
rect 6457 6239 6515 6245
rect 6457 6236 6469 6239
rect 5675 6208 6469 6236
rect 5675 6205 5687 6208
rect 5629 6199 5687 6205
rect 6457 6205 6469 6208
rect 6503 6205 6515 6239
rect 7668 6236 7696 6412
rect 8113 6409 8125 6412
rect 8159 6409 8171 6443
rect 9585 6443 9643 6449
rect 9585 6440 9597 6443
rect 8113 6403 8171 6409
rect 8220 6412 9597 6440
rect 8220 6384 8248 6412
rect 9585 6409 9597 6412
rect 9631 6440 9643 6443
rect 10502 6440 10508 6452
rect 9631 6412 10508 6440
rect 9631 6409 9643 6412
rect 9585 6403 9643 6409
rect 10502 6400 10508 6412
rect 10560 6400 10566 6452
rect 11790 6400 11796 6452
rect 11848 6440 11854 6452
rect 11885 6443 11943 6449
rect 11885 6440 11897 6443
rect 11848 6412 11897 6440
rect 11848 6400 11854 6412
rect 11885 6409 11897 6412
rect 11931 6409 11943 6443
rect 11885 6403 11943 6409
rect 12250 6400 12256 6452
rect 12308 6400 12314 6452
rect 20349 6443 20407 6449
rect 20349 6409 20361 6443
rect 20395 6409 20407 6443
rect 20349 6403 20407 6409
rect 20717 6443 20775 6449
rect 20717 6409 20729 6443
rect 20763 6440 20775 6443
rect 21082 6440 21088 6452
rect 20763 6412 21088 6440
rect 20763 6409 20775 6412
rect 20717 6403 20775 6409
rect 7745 6375 7803 6381
rect 7745 6341 7757 6375
rect 7791 6372 7803 6375
rect 7834 6372 7840 6384
rect 7791 6344 7840 6372
rect 7791 6341 7803 6344
rect 7745 6335 7803 6341
rect 7834 6332 7840 6344
rect 7892 6332 7898 6384
rect 7975 6341 8033 6347
rect 7975 6307 7987 6341
rect 8021 6307 8033 6341
rect 8202 6332 8208 6384
rect 8260 6332 8266 6384
rect 8938 6372 8944 6384
rect 8312 6344 8944 6372
rect 8312 6316 8340 6344
rect 8938 6332 8944 6344
rect 8996 6372 9002 6384
rect 9214 6372 9220 6384
rect 8996 6344 9220 6372
rect 8996 6332 9002 6344
rect 9214 6332 9220 6344
rect 9272 6332 9278 6384
rect 9306 6332 9312 6384
rect 9364 6372 9370 6384
rect 9364 6344 12434 6372
rect 9364 6332 9370 6344
rect 7975 6304 8033 6307
rect 8294 6304 8300 6316
rect 7975 6301 8300 6304
rect 7976 6276 8300 6301
rect 8294 6264 8300 6276
rect 8352 6264 8358 6316
rect 8754 6264 8760 6316
rect 8812 6264 8818 6316
rect 8846 6264 8852 6316
rect 8904 6304 8910 6316
rect 9401 6307 9459 6313
rect 9401 6304 9413 6307
rect 8904 6276 9413 6304
rect 8904 6264 8910 6276
rect 9401 6273 9413 6276
rect 9447 6273 9459 6307
rect 9401 6267 9459 6273
rect 9677 6307 9735 6313
rect 9677 6273 9689 6307
rect 9723 6304 9735 6307
rect 9858 6304 9864 6316
rect 9723 6276 9864 6304
rect 9723 6273 9735 6276
rect 9677 6267 9735 6273
rect 9858 6264 9864 6276
rect 9916 6264 9922 6316
rect 9950 6264 9956 6316
rect 10008 6264 10014 6316
rect 10152 6313 10180 6344
rect 10137 6307 10195 6313
rect 10137 6273 10149 6307
rect 10183 6273 10195 6307
rect 10137 6267 10195 6273
rect 11057 6307 11115 6313
rect 11057 6273 11069 6307
rect 11103 6304 11115 6307
rect 11422 6304 11428 6316
rect 11103 6276 11428 6304
rect 11103 6273 11115 6276
rect 11057 6267 11115 6273
rect 11422 6264 11428 6276
rect 11480 6264 11486 6316
rect 12406 6304 12434 6344
rect 12618 6332 12624 6384
rect 12676 6372 12682 6384
rect 13354 6372 13360 6384
rect 12676 6344 13360 6372
rect 12676 6332 12682 6344
rect 13354 6332 13360 6344
rect 13412 6332 13418 6384
rect 18785 6375 18843 6381
rect 18785 6372 18797 6375
rect 17972 6344 18797 6372
rect 13541 6307 13599 6313
rect 13541 6304 13553 6307
rect 12406 6276 13553 6304
rect 13541 6273 13553 6276
rect 13587 6304 13599 6307
rect 13906 6304 13912 6316
rect 13587 6276 13912 6304
rect 13587 6273 13599 6276
rect 13541 6267 13599 6273
rect 13906 6264 13912 6276
rect 13964 6264 13970 6316
rect 15838 6264 15844 6316
rect 15896 6264 15902 6316
rect 16761 6307 16819 6313
rect 16761 6273 16773 6307
rect 16807 6304 16819 6307
rect 16942 6304 16948 6316
rect 16807 6276 16948 6304
rect 16807 6273 16819 6276
rect 16761 6267 16819 6273
rect 16942 6264 16948 6276
rect 17000 6264 17006 6316
rect 17678 6264 17684 6316
rect 17736 6264 17742 6316
rect 17972 6313 18000 6344
rect 18785 6341 18797 6344
rect 18831 6341 18843 6375
rect 18785 6335 18843 6341
rect 17957 6307 18015 6313
rect 17957 6273 17969 6307
rect 18003 6273 18015 6307
rect 17957 6267 18015 6273
rect 18141 6307 18199 6313
rect 18141 6273 18153 6307
rect 18187 6273 18199 6307
rect 18141 6267 18199 6273
rect 8570 6236 8576 6248
rect 7668 6208 8576 6236
rect 6457 6199 6515 6205
rect 8570 6196 8576 6208
rect 8628 6236 8634 6248
rect 8665 6239 8723 6245
rect 8665 6236 8677 6239
rect 8628 6208 8677 6236
rect 8628 6196 8634 6208
rect 8665 6205 8677 6208
rect 8711 6236 8723 6239
rect 10318 6236 10324 6248
rect 8711 6208 10324 6236
rect 8711 6205 8723 6208
rect 8665 6199 8723 6205
rect 10318 6196 10324 6208
rect 10376 6196 10382 6248
rect 12345 6239 12403 6245
rect 12345 6205 12357 6239
rect 12391 6205 12403 6239
rect 12345 6199 12403 6205
rect 12529 6239 12587 6245
rect 12529 6205 12541 6239
rect 12575 6236 12587 6239
rect 13814 6236 13820 6248
rect 12575 6208 13820 6236
rect 12575 6205 12587 6208
rect 12529 6199 12587 6205
rect 5997 6171 6055 6177
rect 5997 6168 6009 6171
rect 4816 6140 6009 6168
rect 4341 6131 4399 6137
rect 5997 6137 6009 6140
rect 6043 6168 6055 6171
rect 6641 6171 6699 6177
rect 6641 6168 6653 6171
rect 6043 6140 6653 6168
rect 6043 6137 6055 6140
rect 5997 6131 6055 6137
rect 6641 6137 6653 6140
rect 6687 6137 6699 6171
rect 6641 6131 6699 6137
rect 8128 6140 8708 6168
rect 2866 6060 2872 6112
rect 2924 6100 2930 6112
rect 7650 6100 7656 6112
rect 2924 6072 7656 6100
rect 2924 6060 2930 6072
rect 7650 6060 7656 6072
rect 7708 6060 7714 6112
rect 7742 6060 7748 6112
rect 7800 6100 7806 6112
rect 7929 6103 7987 6109
rect 7929 6100 7941 6103
rect 7800 6072 7941 6100
rect 7800 6060 7806 6072
rect 7929 6069 7941 6072
rect 7975 6100 7987 6103
rect 8128 6100 8156 6140
rect 8680 6112 8708 6140
rect 8754 6128 8760 6180
rect 8812 6168 8818 6180
rect 9398 6168 9404 6180
rect 8812 6140 9404 6168
rect 8812 6128 8818 6140
rect 9398 6128 9404 6140
rect 9456 6128 9462 6180
rect 9766 6128 9772 6180
rect 9824 6168 9830 6180
rect 10873 6171 10931 6177
rect 10873 6168 10885 6171
rect 9824 6140 10885 6168
rect 9824 6128 9830 6140
rect 10873 6137 10885 6140
rect 10919 6137 10931 6171
rect 12360 6168 12388 6199
rect 13814 6196 13820 6208
rect 13872 6196 13878 6248
rect 14458 6196 14464 6248
rect 14516 6196 14522 6248
rect 14737 6239 14795 6245
rect 14737 6205 14749 6239
rect 14783 6236 14795 6239
rect 15102 6236 15108 6248
rect 14783 6208 15108 6236
rect 14783 6205 14795 6208
rect 14737 6199 14795 6205
rect 15102 6196 15108 6208
rect 15160 6196 15166 6248
rect 18156 6236 18184 6267
rect 18598 6264 18604 6316
rect 18656 6304 18662 6316
rect 19150 6304 19156 6316
rect 18656 6276 19156 6304
rect 18656 6264 18662 6276
rect 19150 6264 19156 6276
rect 19208 6264 19214 6316
rect 20073 6307 20131 6313
rect 20073 6273 20085 6307
rect 20119 6304 20131 6307
rect 20364 6304 20392 6403
rect 21082 6400 21088 6412
rect 21140 6400 21146 6452
rect 21358 6400 21364 6452
rect 21416 6400 21422 6452
rect 21913 6443 21971 6449
rect 21913 6409 21925 6443
rect 21959 6409 21971 6443
rect 21913 6403 21971 6409
rect 20119 6276 20392 6304
rect 21545 6307 21603 6313
rect 20119 6273 20131 6276
rect 20073 6267 20131 6273
rect 21545 6273 21557 6307
rect 21591 6304 21603 6307
rect 21928 6304 21956 6403
rect 25038 6400 25044 6452
rect 25096 6400 25102 6452
rect 22370 6332 22376 6384
rect 22428 6332 22434 6384
rect 23658 6332 23664 6384
rect 23716 6372 23722 6384
rect 23716 6344 24058 6372
rect 23716 6332 23722 6344
rect 21591 6276 21956 6304
rect 21591 6273 21603 6276
rect 21545 6267 21603 6273
rect 22094 6264 22100 6316
rect 22152 6304 22158 6316
rect 22281 6307 22339 6313
rect 22281 6304 22293 6307
rect 22152 6276 22293 6304
rect 22152 6264 22158 6276
rect 22281 6273 22293 6276
rect 22327 6273 22339 6307
rect 22388 6304 22416 6332
rect 23106 6304 23112 6316
rect 22388 6276 23112 6304
rect 22281 6267 22339 6273
rect 19610 6236 19616 6248
rect 18156 6208 19616 6236
rect 19610 6196 19616 6208
rect 19668 6196 19674 6248
rect 20622 6196 20628 6248
rect 20680 6236 20686 6248
rect 20809 6239 20867 6245
rect 20809 6236 20821 6239
rect 20680 6208 20821 6236
rect 20680 6196 20686 6208
rect 20809 6205 20821 6208
rect 20855 6205 20867 6239
rect 20809 6199 20867 6205
rect 20898 6196 20904 6248
rect 20956 6196 20962 6248
rect 22296 6168 22324 6267
rect 23106 6264 23112 6276
rect 23164 6304 23170 6316
rect 23293 6307 23351 6313
rect 23293 6304 23305 6307
rect 23164 6276 23305 6304
rect 23164 6264 23170 6276
rect 23293 6273 23305 6276
rect 23339 6273 23351 6307
rect 23293 6267 23351 6273
rect 22370 6196 22376 6248
rect 22428 6196 22434 6248
rect 22557 6239 22615 6245
rect 22557 6205 22569 6239
rect 22603 6236 22615 6239
rect 22646 6236 22652 6248
rect 22603 6208 22652 6236
rect 22603 6205 22615 6208
rect 22557 6199 22615 6205
rect 22646 6196 22652 6208
rect 22704 6196 22710 6248
rect 23569 6239 23627 6245
rect 23569 6205 23581 6239
rect 23615 6236 23627 6239
rect 23934 6236 23940 6248
rect 23615 6208 23940 6236
rect 23615 6205 23627 6208
rect 23569 6199 23627 6205
rect 23934 6196 23940 6208
rect 23992 6196 23998 6248
rect 12360 6140 14596 6168
rect 10873 6131 10931 6137
rect 7975 6072 8156 6100
rect 7975 6069 7987 6072
rect 7929 6063 7987 6069
rect 8202 6060 8208 6112
rect 8260 6100 8266 6112
rect 8389 6103 8447 6109
rect 8389 6100 8401 6103
rect 8260 6072 8401 6100
rect 8260 6060 8266 6072
rect 8389 6069 8401 6072
rect 8435 6069 8447 6103
rect 8389 6063 8447 6069
rect 8662 6060 8668 6112
rect 8720 6060 8726 6112
rect 9217 6103 9275 6109
rect 9217 6069 9229 6103
rect 9263 6100 9275 6103
rect 9582 6100 9588 6112
rect 9263 6072 9588 6100
rect 9263 6069 9275 6072
rect 9217 6063 9275 6069
rect 9582 6060 9588 6072
rect 9640 6060 9646 6112
rect 10042 6060 10048 6112
rect 10100 6100 10106 6112
rect 10137 6103 10195 6109
rect 10137 6100 10149 6103
rect 10100 6072 10149 6100
rect 10100 6060 10106 6072
rect 10137 6069 10149 6072
rect 10183 6069 10195 6103
rect 14568 6100 14596 6140
rect 15764 6140 22324 6168
rect 15764 6100 15792 6140
rect 14568 6072 15792 6100
rect 10137 6063 10195 6069
rect 15930 6060 15936 6112
rect 15988 6100 15994 6112
rect 16209 6103 16267 6109
rect 16209 6100 16221 6103
rect 15988 6072 16221 6100
rect 15988 6060 15994 6072
rect 16209 6069 16221 6072
rect 16255 6069 16267 6103
rect 16209 6063 16267 6069
rect 16945 6103 17003 6109
rect 16945 6069 16957 6103
rect 16991 6100 17003 6103
rect 17034 6100 17040 6112
rect 16991 6072 17040 6100
rect 16991 6069 17003 6072
rect 16945 6063 17003 6069
rect 17034 6060 17040 6072
rect 17092 6060 17098 6112
rect 17218 6060 17224 6112
rect 17276 6100 17282 6112
rect 17497 6103 17555 6109
rect 17497 6100 17509 6103
rect 17276 6072 17509 6100
rect 17276 6060 17282 6072
rect 17497 6069 17509 6072
rect 17543 6069 17555 6103
rect 17497 6063 17555 6069
rect 18141 6103 18199 6109
rect 18141 6069 18153 6103
rect 18187 6100 18199 6103
rect 18230 6100 18236 6112
rect 18187 6072 18236 6100
rect 18187 6069 18199 6072
rect 18141 6063 18199 6069
rect 18230 6060 18236 6072
rect 18288 6060 18294 6112
rect 18693 6103 18751 6109
rect 18693 6069 18705 6103
rect 18739 6100 18751 6103
rect 19702 6100 19708 6112
rect 18739 6072 19708 6100
rect 18739 6069 18751 6072
rect 18693 6063 18751 6069
rect 19702 6060 19708 6072
rect 19760 6060 19766 6112
rect 19794 6060 19800 6112
rect 19852 6100 19858 6112
rect 19889 6103 19947 6109
rect 19889 6100 19901 6103
rect 19852 6072 19901 6100
rect 19852 6060 19858 6072
rect 19889 6069 19901 6072
rect 19935 6069 19947 6103
rect 19889 6063 19947 6069
rect 1104 6010 25852 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 12214 6010
rect 12266 5958 12278 6010
rect 12330 5958 12342 6010
rect 12394 5958 12406 6010
rect 12458 5958 12470 6010
rect 12522 5958 20214 6010
rect 20266 5958 20278 6010
rect 20330 5958 20342 6010
rect 20394 5958 20406 6010
rect 20458 5958 20470 6010
rect 20522 5958 25852 6010
rect 1104 5936 25852 5958
rect 4540 5868 5120 5896
rect 2774 5788 2780 5840
rect 2832 5788 2838 5840
rect 4540 5769 4568 5868
rect 4706 5828 4712 5840
rect 4632 5800 4712 5828
rect 4632 5769 4660 5800
rect 4706 5788 4712 5800
rect 4764 5788 4770 5840
rect 5092 5828 5120 5868
rect 5166 5856 5172 5908
rect 5224 5896 5230 5908
rect 5353 5899 5411 5905
rect 5353 5896 5365 5899
rect 5224 5868 5365 5896
rect 5224 5856 5230 5868
rect 5353 5865 5365 5868
rect 5399 5865 5411 5899
rect 5353 5859 5411 5865
rect 6196 5868 7052 5896
rect 6196 5828 6224 5868
rect 5092 5800 6224 5828
rect 6273 5831 6331 5837
rect 6273 5797 6285 5831
rect 6319 5828 6331 5831
rect 6914 5828 6920 5840
rect 6319 5800 6920 5828
rect 6319 5797 6331 5800
rect 6273 5791 6331 5797
rect 4525 5763 4583 5769
rect 4525 5729 4537 5763
rect 4571 5729 4583 5763
rect 4525 5723 4583 5729
rect 4617 5763 4675 5769
rect 4617 5729 4629 5763
rect 4663 5729 4675 5763
rect 5813 5763 5871 5769
rect 5813 5760 5825 5763
rect 4617 5723 4675 5729
rect 5276 5732 5825 5760
rect 5276 5704 5304 5732
rect 5813 5729 5825 5732
rect 5859 5729 5871 5763
rect 5813 5723 5871 5729
rect 2225 5695 2283 5701
rect 2225 5661 2237 5695
rect 2271 5661 2283 5695
rect 2225 5655 2283 5661
rect 2240 5624 2268 5655
rect 2498 5652 2504 5704
rect 2556 5692 2562 5704
rect 2593 5695 2651 5701
rect 2593 5692 2605 5695
rect 2556 5664 2605 5692
rect 2556 5652 2562 5664
rect 2593 5661 2605 5664
rect 2639 5661 2651 5695
rect 2593 5655 2651 5661
rect 2777 5695 2835 5701
rect 2777 5661 2789 5695
rect 2823 5692 2835 5695
rect 2866 5692 2872 5704
rect 2823 5664 2872 5692
rect 2823 5661 2835 5664
rect 2777 5655 2835 5661
rect 2866 5652 2872 5664
rect 2924 5652 2930 5704
rect 3326 5652 3332 5704
rect 3384 5701 3390 5704
rect 3510 5701 3516 5704
rect 3384 5695 3417 5701
rect 3405 5661 3417 5695
rect 3384 5655 3417 5661
rect 3506 5655 3516 5701
rect 3384 5652 3390 5655
rect 3510 5652 3516 5655
rect 3568 5652 3574 5704
rect 4706 5652 4712 5704
rect 4764 5652 4770 5704
rect 4801 5695 4859 5701
rect 4801 5661 4813 5695
rect 4847 5692 4859 5695
rect 5166 5692 5172 5704
rect 4847 5664 5172 5692
rect 4847 5661 4859 5664
rect 4801 5655 4859 5661
rect 5166 5652 5172 5664
rect 5224 5652 5230 5704
rect 5258 5652 5264 5704
rect 5316 5652 5322 5704
rect 5445 5695 5503 5701
rect 5445 5661 5457 5695
rect 5491 5692 5503 5695
rect 5905 5695 5963 5701
rect 5905 5692 5917 5695
rect 5491 5664 5917 5692
rect 5491 5661 5503 5664
rect 5445 5655 5503 5661
rect 5905 5661 5917 5664
rect 5951 5692 5963 5695
rect 6086 5692 6092 5704
rect 5951 5664 6092 5692
rect 5951 5661 5963 5664
rect 5905 5655 5963 5661
rect 6086 5652 6092 5664
rect 6144 5652 6150 5704
rect 6288 5692 6316 5791
rect 6914 5788 6920 5800
rect 6972 5788 6978 5840
rect 7024 5828 7052 5868
rect 7098 5856 7104 5908
rect 7156 5856 7162 5908
rect 11422 5896 11428 5908
rect 7576 5868 11428 5896
rect 7576 5828 7604 5868
rect 11422 5856 11428 5868
rect 11480 5856 11486 5908
rect 11517 5899 11575 5905
rect 11517 5865 11529 5899
rect 11563 5896 11575 5899
rect 12066 5896 12072 5908
rect 11563 5868 12072 5896
rect 11563 5865 11575 5868
rect 11517 5859 11575 5865
rect 12066 5856 12072 5868
rect 12124 5856 12130 5908
rect 12176 5868 13768 5896
rect 7024 5800 7604 5828
rect 7653 5831 7711 5837
rect 7653 5797 7665 5831
rect 7699 5828 7711 5831
rect 8938 5828 8944 5840
rect 7699 5800 8944 5828
rect 7699 5797 7711 5800
rect 7653 5791 7711 5797
rect 8938 5788 8944 5800
rect 8996 5788 9002 5840
rect 12176 5828 12204 5868
rect 13740 5840 13768 5868
rect 15102 5856 15108 5908
rect 15160 5856 15166 5908
rect 19426 5896 19432 5908
rect 15212 5868 19432 5896
rect 10428 5800 12204 5828
rect 13541 5831 13599 5837
rect 8294 5760 8300 5772
rect 7944 5732 8300 5760
rect 6549 5695 6607 5701
rect 6549 5692 6561 5695
rect 6288 5664 6561 5692
rect 6549 5661 6561 5664
rect 6595 5661 6607 5695
rect 6549 5655 6607 5661
rect 6825 5695 6883 5701
rect 6825 5661 6837 5695
rect 6871 5692 6883 5695
rect 6871 5664 7328 5692
rect 6871 5661 6883 5664
rect 6825 5655 6883 5661
rect 3234 5624 3240 5636
rect 2240 5596 3240 5624
rect 3234 5584 3240 5596
rect 3292 5584 3298 5636
rect 5994 5584 6000 5636
rect 6052 5624 6058 5636
rect 6641 5627 6699 5633
rect 6052 5596 6408 5624
rect 6052 5584 6058 5596
rect 2038 5516 2044 5568
rect 2096 5516 2102 5568
rect 3142 5516 3148 5568
rect 3200 5516 3206 5568
rect 4985 5559 5043 5565
rect 4985 5525 4997 5559
rect 5031 5556 5043 5559
rect 5902 5556 5908 5568
rect 5031 5528 5908 5556
rect 5031 5525 5043 5528
rect 4985 5519 5043 5525
rect 5902 5516 5908 5528
rect 5960 5516 5966 5568
rect 6380 5556 6408 5596
rect 6641 5593 6653 5627
rect 6687 5624 6699 5627
rect 7006 5624 7012 5636
rect 6687 5596 7012 5624
rect 6687 5593 6699 5596
rect 6641 5587 6699 5593
rect 7006 5584 7012 5596
rect 7064 5584 7070 5636
rect 7098 5584 7104 5636
rect 7156 5584 7162 5636
rect 7300 5624 7328 5664
rect 7374 5652 7380 5704
rect 7432 5652 7438 5704
rect 7653 5695 7711 5701
rect 7653 5661 7665 5695
rect 7699 5692 7711 5695
rect 7834 5692 7840 5704
rect 7699 5664 7840 5692
rect 7699 5661 7711 5664
rect 7653 5655 7711 5661
rect 7834 5652 7840 5664
rect 7892 5652 7898 5704
rect 7944 5701 7972 5732
rect 8294 5720 8300 5732
rect 8352 5720 8358 5772
rect 10428 5760 10456 5800
rect 13541 5797 13553 5831
rect 13587 5828 13599 5831
rect 13630 5828 13636 5840
rect 13587 5800 13636 5828
rect 13587 5797 13599 5800
rect 13541 5791 13599 5797
rect 13630 5788 13636 5800
rect 13688 5788 13694 5840
rect 13722 5788 13728 5840
rect 13780 5828 13786 5840
rect 15212 5828 15240 5868
rect 19426 5856 19432 5868
rect 19484 5856 19490 5908
rect 23658 5856 23664 5908
rect 23716 5856 23722 5908
rect 13780 5800 15240 5828
rect 15565 5831 15623 5837
rect 13780 5788 13786 5800
rect 15565 5797 15577 5831
rect 15611 5797 15623 5831
rect 15565 5791 15623 5797
rect 8404 5732 10456 5760
rect 12897 5763 12955 5769
rect 7929 5695 7987 5701
rect 7929 5661 7941 5695
rect 7975 5661 7987 5695
rect 7929 5655 7987 5661
rect 8202 5652 8208 5704
rect 8260 5652 8266 5704
rect 7558 5624 7564 5636
rect 7300 5596 7564 5624
rect 7558 5584 7564 5596
rect 7616 5584 7622 5636
rect 7668 5596 7972 5624
rect 7668 5568 7696 5596
rect 6733 5559 6791 5565
rect 6733 5556 6745 5559
rect 6380 5528 6745 5556
rect 6733 5525 6745 5528
rect 6779 5556 6791 5559
rect 7285 5559 7343 5565
rect 7285 5556 7297 5559
rect 6779 5528 7297 5556
rect 6779 5525 6791 5528
rect 6733 5519 6791 5525
rect 7285 5525 7297 5528
rect 7331 5525 7343 5559
rect 7285 5519 7343 5525
rect 7650 5516 7656 5568
rect 7708 5516 7714 5568
rect 7742 5516 7748 5568
rect 7800 5556 7806 5568
rect 7837 5559 7895 5565
rect 7837 5556 7849 5559
rect 7800 5528 7849 5556
rect 7800 5516 7806 5528
rect 7837 5525 7849 5528
rect 7883 5525 7895 5559
rect 7944 5556 7972 5596
rect 8018 5584 8024 5636
rect 8076 5624 8082 5636
rect 8297 5627 8355 5633
rect 8297 5624 8309 5627
rect 8076 5596 8309 5624
rect 8076 5584 8082 5596
rect 8297 5593 8309 5596
rect 8343 5593 8355 5627
rect 8297 5587 8355 5593
rect 8404 5556 8432 5732
rect 12897 5729 12909 5763
rect 12943 5760 12955 5763
rect 13262 5760 13268 5772
rect 12943 5732 13268 5760
rect 12943 5729 12955 5732
rect 12897 5723 12955 5729
rect 13262 5720 13268 5732
rect 13320 5760 13326 5772
rect 13814 5760 13820 5772
rect 13320 5732 13820 5760
rect 13320 5720 13326 5732
rect 13814 5720 13820 5732
rect 13872 5720 13878 5772
rect 8481 5695 8539 5701
rect 8481 5661 8493 5695
rect 8527 5692 8539 5695
rect 8754 5692 8760 5704
rect 8527 5664 8760 5692
rect 8527 5661 8539 5664
rect 8481 5655 8539 5661
rect 8754 5652 8760 5664
rect 8812 5652 8818 5704
rect 9030 5652 9036 5704
rect 9088 5652 9094 5704
rect 11333 5695 11391 5701
rect 11333 5661 11345 5695
rect 11379 5692 11391 5695
rect 11422 5692 11428 5704
rect 11379 5664 11428 5692
rect 11379 5661 11391 5664
rect 11333 5655 11391 5661
rect 11422 5652 11428 5664
rect 11480 5652 11486 5704
rect 12713 5695 12771 5701
rect 12713 5661 12725 5695
rect 12759 5692 12771 5695
rect 15289 5695 15347 5701
rect 12759 5664 14412 5692
rect 12759 5661 12771 5664
rect 12713 5655 12771 5661
rect 8665 5627 8723 5633
rect 8665 5593 8677 5627
rect 8711 5624 8723 5627
rect 9309 5627 9367 5633
rect 9309 5624 9321 5627
rect 8711 5596 9321 5624
rect 8711 5593 8723 5596
rect 8665 5587 8723 5593
rect 9309 5593 9321 5596
rect 9355 5593 9367 5627
rect 9309 5587 9367 5593
rect 10042 5584 10048 5636
rect 10100 5584 10106 5636
rect 11974 5584 11980 5636
rect 12032 5624 12038 5636
rect 12621 5627 12679 5633
rect 12621 5624 12633 5627
rect 12032 5596 12633 5624
rect 12032 5584 12038 5596
rect 12621 5593 12633 5596
rect 12667 5593 12679 5627
rect 12621 5587 12679 5593
rect 13354 5584 13360 5636
rect 13412 5584 13418 5636
rect 7944 5528 8432 5556
rect 7837 5519 7895 5525
rect 9490 5516 9496 5568
rect 9548 5556 9554 5568
rect 10781 5559 10839 5565
rect 10781 5556 10793 5559
rect 9548 5528 10793 5556
rect 9548 5516 9554 5528
rect 10781 5525 10793 5528
rect 10827 5525 10839 5559
rect 10781 5519 10839 5525
rect 11514 5516 11520 5568
rect 11572 5516 11578 5568
rect 12066 5516 12072 5568
rect 12124 5556 12130 5568
rect 12253 5559 12311 5565
rect 12253 5556 12265 5559
rect 12124 5528 12265 5556
rect 12124 5516 12130 5528
rect 12253 5525 12265 5528
rect 12299 5525 12311 5559
rect 14384 5556 14412 5664
rect 15289 5661 15301 5695
rect 15335 5692 15347 5695
rect 15580 5692 15608 5791
rect 16114 5720 16120 5772
rect 16172 5720 16178 5772
rect 19518 5760 19524 5772
rect 16960 5732 19524 5760
rect 16960 5701 16988 5732
rect 19518 5720 19524 5732
rect 19576 5720 19582 5772
rect 19794 5720 19800 5772
rect 19852 5720 19858 5772
rect 16945 5695 17003 5701
rect 16945 5692 16957 5695
rect 15335 5664 15608 5692
rect 16684 5664 16957 5692
rect 15335 5661 15347 5664
rect 15289 5655 15347 5661
rect 16684 5636 16712 5664
rect 16945 5661 16957 5664
rect 16991 5661 17003 5695
rect 16945 5655 17003 5661
rect 23382 5652 23388 5704
rect 23440 5652 23446 5704
rect 23566 5652 23572 5704
rect 23624 5692 23630 5704
rect 23661 5695 23719 5701
rect 23661 5692 23673 5695
rect 23624 5664 23673 5692
rect 23624 5652 23630 5664
rect 23661 5661 23673 5664
rect 23707 5661 23719 5695
rect 23661 5655 23719 5661
rect 23750 5652 23756 5704
rect 23808 5692 23814 5704
rect 23845 5695 23903 5701
rect 23845 5692 23857 5695
rect 23808 5664 23857 5692
rect 23808 5652 23814 5664
rect 23845 5661 23857 5664
rect 23891 5661 23903 5695
rect 23845 5655 23903 5661
rect 14458 5584 14464 5636
rect 14516 5624 14522 5636
rect 16666 5624 16672 5636
rect 14516 5596 16672 5624
rect 14516 5584 14522 5596
rect 16666 5584 16672 5596
rect 16724 5584 16730 5636
rect 17218 5584 17224 5636
rect 17276 5584 17282 5636
rect 18230 5584 18236 5636
rect 18288 5584 18294 5636
rect 20806 5584 20812 5636
rect 20864 5584 20870 5636
rect 15930 5556 15936 5568
rect 14384 5528 15936 5556
rect 12253 5519 12311 5525
rect 15930 5516 15936 5528
rect 15988 5516 15994 5568
rect 16025 5559 16083 5565
rect 16025 5525 16037 5559
rect 16071 5556 16083 5559
rect 18138 5556 18144 5568
rect 16071 5528 18144 5556
rect 16071 5525 16083 5528
rect 16025 5519 16083 5525
rect 18138 5516 18144 5528
rect 18196 5556 18202 5568
rect 18693 5559 18751 5565
rect 18693 5556 18705 5559
rect 18196 5528 18705 5556
rect 18196 5516 18202 5528
rect 18693 5525 18705 5528
rect 18739 5525 18751 5559
rect 18693 5519 18751 5525
rect 20162 5516 20168 5568
rect 20220 5556 20226 5568
rect 20622 5556 20628 5568
rect 20220 5528 20628 5556
rect 20220 5516 20226 5528
rect 20622 5516 20628 5528
rect 20680 5556 20686 5568
rect 21269 5559 21327 5565
rect 21269 5556 21281 5559
rect 20680 5528 21281 5556
rect 20680 5516 20686 5528
rect 21269 5525 21281 5528
rect 21315 5525 21327 5559
rect 21269 5519 21327 5525
rect 23201 5559 23259 5565
rect 23201 5525 23213 5559
rect 23247 5556 23259 5559
rect 23290 5556 23296 5568
rect 23247 5528 23296 5556
rect 23247 5525 23259 5528
rect 23201 5519 23259 5525
rect 23290 5516 23296 5528
rect 23348 5516 23354 5568
rect 1104 5466 25852 5488
rect 1104 5414 8214 5466
rect 8266 5414 8278 5466
rect 8330 5414 8342 5466
rect 8394 5414 8406 5466
rect 8458 5414 8470 5466
rect 8522 5414 16214 5466
rect 16266 5414 16278 5466
rect 16330 5414 16342 5466
rect 16394 5414 16406 5466
rect 16458 5414 16470 5466
rect 16522 5414 24214 5466
rect 24266 5414 24278 5466
rect 24330 5414 24342 5466
rect 24394 5414 24406 5466
rect 24458 5414 24470 5466
rect 24522 5414 25852 5466
rect 1104 5392 25852 5414
rect 3234 5312 3240 5364
rect 3292 5352 3298 5364
rect 3513 5355 3571 5361
rect 3513 5352 3525 5355
rect 3292 5324 3525 5352
rect 3292 5312 3298 5324
rect 3513 5321 3525 5324
rect 3559 5321 3571 5355
rect 3513 5315 3571 5321
rect 3602 5312 3608 5364
rect 3660 5352 3666 5364
rect 3881 5355 3939 5361
rect 3881 5352 3893 5355
rect 3660 5324 3893 5352
rect 3660 5312 3666 5324
rect 3881 5321 3893 5324
rect 3927 5321 3939 5355
rect 3881 5315 3939 5321
rect 3973 5355 4031 5361
rect 3973 5321 3985 5355
rect 4019 5352 4031 5355
rect 6457 5355 6515 5361
rect 6457 5352 6469 5355
rect 4019 5324 6469 5352
rect 4019 5321 4031 5324
rect 3973 5315 4031 5321
rect 6457 5321 6469 5324
rect 6503 5321 6515 5355
rect 6457 5315 6515 5321
rect 7006 5312 7012 5364
rect 7064 5352 7070 5364
rect 7469 5355 7527 5361
rect 7469 5352 7481 5355
rect 7064 5324 7481 5352
rect 7064 5312 7070 5324
rect 7469 5321 7481 5324
rect 7515 5352 7527 5355
rect 7650 5352 7656 5364
rect 7515 5324 7656 5352
rect 7515 5321 7527 5324
rect 7469 5315 7527 5321
rect 7650 5312 7656 5324
rect 7708 5312 7714 5364
rect 7834 5312 7840 5364
rect 7892 5352 7898 5364
rect 8113 5355 8171 5361
rect 8113 5352 8125 5355
rect 7892 5324 8125 5352
rect 7892 5312 7898 5324
rect 8113 5321 8125 5324
rect 8159 5321 8171 5355
rect 8113 5315 8171 5321
rect 8938 5312 8944 5364
rect 8996 5352 9002 5364
rect 8996 5324 9720 5352
rect 8996 5312 9002 5324
rect 1765 5287 1823 5293
rect 1765 5253 1777 5287
rect 1811 5284 1823 5287
rect 2038 5284 2044 5296
rect 1811 5256 2044 5284
rect 1811 5253 1823 5256
rect 1765 5247 1823 5253
rect 2038 5244 2044 5256
rect 2096 5244 2102 5296
rect 2774 5244 2780 5296
rect 2832 5244 2838 5296
rect 3786 5244 3792 5296
rect 3844 5284 3850 5296
rect 4798 5284 4804 5296
rect 3844 5256 4804 5284
rect 3844 5244 3850 5256
rect 4798 5244 4804 5256
rect 4856 5244 4862 5296
rect 5721 5287 5779 5293
rect 5721 5253 5733 5287
rect 5767 5284 5779 5287
rect 5767 5256 6868 5284
rect 5767 5253 5779 5256
rect 5721 5247 5779 5253
rect 1486 5176 1492 5228
rect 1544 5176 1550 5228
rect 3326 5176 3332 5228
rect 3384 5216 3390 5228
rect 3384 5188 4476 5216
rect 3384 5176 3390 5188
rect 3237 5151 3295 5157
rect 3237 5117 3249 5151
rect 3283 5148 3295 5151
rect 3510 5148 3516 5160
rect 3283 5120 3516 5148
rect 3283 5117 3295 5120
rect 3237 5111 3295 5117
rect 3510 5108 3516 5120
rect 3568 5108 3574 5160
rect 3970 5108 3976 5160
rect 4028 5148 4034 5160
rect 4065 5151 4123 5157
rect 4065 5148 4077 5151
rect 4028 5120 4077 5148
rect 4028 5108 4034 5120
rect 4065 5117 4077 5120
rect 4111 5117 4123 5151
rect 4448 5148 4476 5188
rect 4522 5176 4528 5228
rect 4580 5176 4586 5228
rect 4706 5225 4712 5228
rect 4673 5219 4712 5225
rect 4673 5185 4685 5219
rect 4673 5179 4712 5185
rect 4706 5176 4712 5179
rect 4764 5176 4770 5228
rect 4890 5176 4896 5228
rect 4948 5176 4954 5228
rect 4982 5176 4988 5228
rect 5040 5225 5046 5228
rect 5040 5219 5067 5225
rect 5055 5185 5067 5219
rect 5994 5216 6000 5228
rect 5955 5188 6000 5216
rect 5040 5179 5067 5185
rect 5040 5176 5046 5179
rect 5994 5176 6000 5188
rect 6052 5176 6058 5228
rect 6840 5225 6868 5256
rect 6914 5244 6920 5296
rect 6972 5284 6978 5296
rect 7285 5287 7343 5293
rect 7285 5284 7297 5287
rect 6972 5256 7297 5284
rect 6972 5244 6978 5256
rect 7285 5253 7297 5256
rect 7331 5253 7343 5287
rect 7285 5247 7343 5253
rect 9122 5244 9128 5296
rect 9180 5244 9186 5296
rect 9582 5244 9588 5296
rect 9640 5244 9646 5296
rect 9692 5284 9720 5324
rect 9858 5312 9864 5364
rect 9916 5352 9922 5364
rect 10229 5355 10287 5361
rect 10229 5352 10241 5355
rect 9916 5324 10241 5352
rect 9916 5312 9922 5324
rect 10229 5321 10241 5324
rect 10275 5321 10287 5355
rect 10229 5315 10287 5321
rect 14918 5312 14924 5364
rect 14976 5352 14982 5364
rect 15197 5355 15255 5361
rect 15197 5352 15209 5355
rect 14976 5324 15209 5352
rect 14976 5312 14982 5324
rect 15197 5321 15209 5324
rect 15243 5321 15255 5355
rect 15197 5315 15255 5321
rect 15746 5312 15752 5364
rect 15804 5312 15810 5364
rect 16114 5352 16120 5364
rect 15948 5324 16120 5352
rect 9692 5256 10180 5284
rect 6089 5219 6147 5225
rect 6089 5185 6101 5219
rect 6135 5185 6147 5219
rect 6089 5179 6147 5185
rect 6825 5219 6883 5225
rect 6825 5185 6837 5219
rect 6871 5185 6883 5219
rect 6825 5179 6883 5185
rect 5000 5148 5028 5176
rect 4448 5120 5028 5148
rect 4065 5111 4123 5117
rect 5074 5040 5080 5092
rect 5132 5080 5138 5092
rect 5169 5083 5227 5089
rect 5169 5080 5181 5083
rect 5132 5052 5181 5080
rect 5132 5040 5138 5052
rect 5169 5049 5181 5052
rect 5215 5049 5227 5083
rect 6104 5080 6132 5179
rect 7558 5176 7564 5228
rect 7616 5216 7622 5228
rect 7926 5216 7932 5228
rect 7616 5188 7932 5216
rect 7616 5176 7622 5188
rect 7926 5176 7932 5188
rect 7984 5176 7990 5228
rect 10152 5225 10180 5256
rect 12618 5244 12624 5296
rect 12676 5244 12682 5296
rect 13354 5244 13360 5296
rect 13412 5284 13418 5296
rect 13817 5287 13875 5293
rect 13817 5284 13829 5287
rect 13412 5256 13829 5284
rect 13412 5244 13418 5256
rect 13817 5253 13829 5256
rect 13863 5253 13875 5287
rect 15470 5284 15476 5296
rect 13817 5247 13875 5253
rect 14292 5256 15476 5284
rect 10137 5219 10195 5225
rect 10137 5185 10149 5219
rect 10183 5185 10195 5219
rect 10137 5179 10195 5185
rect 10318 5176 10324 5228
rect 10376 5176 10382 5228
rect 10962 5176 10968 5228
rect 11020 5216 11026 5228
rect 11609 5219 11667 5225
rect 11609 5216 11621 5219
rect 11020 5188 11621 5216
rect 11020 5176 11026 5188
rect 11609 5185 11621 5188
rect 11655 5185 11667 5219
rect 11609 5179 11667 5185
rect 13722 5176 13728 5228
rect 13780 5216 13786 5228
rect 14292 5225 14320 5256
rect 15470 5244 15476 5256
rect 15528 5244 15534 5296
rect 14277 5219 14335 5225
rect 14277 5216 14289 5219
rect 13780 5188 14289 5216
rect 13780 5176 13786 5188
rect 14277 5185 14289 5188
rect 14323 5185 14335 5219
rect 14277 5179 14335 5185
rect 14461 5219 14519 5225
rect 14461 5185 14473 5219
rect 14507 5216 14519 5219
rect 14507 5188 14872 5216
rect 14507 5185 14519 5188
rect 14461 5179 14519 5185
rect 6733 5151 6791 5157
rect 6733 5117 6745 5151
rect 6779 5148 6791 5151
rect 7374 5148 7380 5160
rect 6779 5120 7380 5148
rect 6779 5117 6791 5120
rect 6733 5111 6791 5117
rect 7374 5108 7380 5120
rect 7432 5108 7438 5160
rect 9861 5151 9919 5157
rect 9861 5117 9873 5151
rect 9907 5148 9919 5151
rect 10980 5148 11008 5176
rect 9907 5120 11008 5148
rect 9907 5117 9919 5120
rect 9861 5111 9919 5117
rect 11882 5108 11888 5160
rect 11940 5108 11946 5160
rect 7098 5080 7104 5092
rect 6104 5052 7104 5080
rect 5169 5043 5227 5049
rect 7098 5040 7104 5052
rect 7156 5080 7162 5092
rect 7285 5083 7343 5089
rect 7285 5080 7297 5083
rect 7156 5052 7297 5080
rect 7156 5040 7162 5052
rect 7285 5049 7297 5052
rect 7331 5049 7343 5083
rect 7285 5043 7343 5049
rect 14182 5040 14188 5092
rect 14240 5080 14246 5092
rect 14737 5083 14795 5089
rect 14737 5080 14749 5083
rect 14240 5052 14749 5080
rect 14240 5040 14246 5052
rect 14737 5049 14749 5052
rect 14783 5049 14795 5083
rect 14844 5080 14872 5188
rect 15102 5176 15108 5228
rect 15160 5176 15166 5228
rect 15948 5216 15976 5324
rect 16114 5312 16120 5324
rect 16172 5352 16178 5364
rect 16945 5355 17003 5361
rect 16945 5352 16957 5355
rect 16172 5324 16957 5352
rect 16172 5312 16178 5324
rect 16945 5321 16957 5324
rect 16991 5321 17003 5355
rect 16945 5315 17003 5321
rect 17678 5312 17684 5364
rect 17736 5352 17742 5364
rect 17865 5355 17923 5361
rect 17865 5352 17877 5355
rect 17736 5324 17877 5352
rect 17736 5312 17742 5324
rect 17865 5321 17877 5324
rect 17911 5321 17923 5355
rect 17865 5315 17923 5321
rect 18138 5312 18144 5364
rect 18196 5352 18202 5364
rect 18233 5355 18291 5361
rect 18233 5352 18245 5355
rect 18196 5324 18245 5352
rect 18196 5312 18202 5324
rect 18233 5321 18245 5324
rect 18279 5321 18291 5355
rect 18233 5315 18291 5321
rect 18325 5355 18383 5361
rect 18325 5321 18337 5355
rect 18371 5352 18383 5355
rect 20162 5352 20168 5364
rect 18371 5324 20168 5352
rect 18371 5321 18383 5324
rect 18325 5315 18383 5321
rect 20162 5312 20168 5324
rect 20220 5312 20226 5364
rect 20441 5355 20499 5361
rect 20441 5321 20453 5355
rect 20487 5352 20499 5355
rect 20806 5352 20812 5364
rect 20487 5324 20812 5352
rect 20487 5321 20499 5324
rect 20441 5315 20499 5321
rect 20806 5312 20812 5324
rect 20864 5312 20870 5364
rect 21913 5355 21971 5361
rect 21913 5321 21925 5355
rect 21959 5321 21971 5355
rect 21913 5315 21971 5321
rect 22281 5355 22339 5361
rect 22281 5321 22293 5355
rect 22327 5352 22339 5355
rect 22370 5352 22376 5364
rect 22327 5324 22376 5352
rect 22327 5321 22339 5324
rect 22281 5315 22339 5321
rect 19702 5244 19708 5296
rect 19760 5284 19766 5296
rect 19760 5256 20392 5284
rect 19760 5244 19766 5256
rect 15304 5188 15976 5216
rect 14918 5108 14924 5160
rect 14976 5148 14982 5160
rect 15304 5148 15332 5188
rect 16022 5176 16028 5228
rect 16080 5176 16086 5228
rect 16114 5176 16120 5228
rect 16172 5176 16178 5228
rect 16761 5219 16819 5225
rect 16761 5185 16773 5219
rect 16807 5216 16819 5219
rect 16942 5216 16948 5228
rect 16807 5188 16948 5216
rect 16807 5185 16819 5188
rect 16761 5179 16819 5185
rect 16942 5176 16948 5188
rect 17000 5176 17006 5228
rect 19150 5176 19156 5228
rect 19208 5176 19214 5228
rect 19978 5216 19984 5228
rect 19260 5188 19984 5216
rect 14976 5120 15332 5148
rect 15381 5151 15439 5157
rect 14976 5108 14982 5120
rect 15381 5117 15393 5151
rect 15427 5148 15439 5151
rect 17034 5148 17040 5160
rect 15427 5120 17040 5148
rect 15427 5117 15439 5120
rect 15381 5111 15439 5117
rect 17034 5108 17040 5120
rect 17092 5148 17098 5160
rect 18509 5151 18567 5157
rect 18509 5148 18521 5151
rect 17092 5120 18521 5148
rect 17092 5108 17098 5120
rect 18509 5117 18521 5120
rect 18555 5148 18567 5151
rect 19260 5148 19288 5188
rect 19978 5176 19984 5188
rect 20036 5176 20042 5228
rect 20364 5225 20392 5256
rect 20349 5219 20407 5225
rect 20349 5185 20361 5219
rect 20395 5185 20407 5219
rect 20349 5179 20407 5185
rect 20533 5219 20591 5225
rect 20533 5185 20545 5219
rect 20579 5216 20591 5219
rect 20622 5216 20628 5228
rect 20579 5188 20628 5216
rect 20579 5185 20591 5188
rect 20533 5179 20591 5185
rect 20622 5176 20628 5188
rect 20680 5176 20686 5228
rect 21361 5219 21419 5225
rect 21361 5185 21373 5219
rect 21407 5216 21419 5219
rect 21928 5216 21956 5315
rect 22370 5312 22376 5324
rect 22428 5312 22434 5364
rect 23658 5244 23664 5296
rect 23716 5284 23722 5296
rect 23716 5256 23874 5284
rect 23716 5244 23722 5256
rect 21407 5188 21956 5216
rect 22020 5188 22600 5216
rect 21407 5185 21419 5188
rect 21361 5179 21419 5185
rect 18555 5120 19288 5148
rect 19429 5151 19487 5157
rect 18555 5117 18567 5120
rect 18509 5111 18567 5117
rect 19429 5117 19441 5151
rect 19475 5148 19487 5151
rect 20070 5148 20076 5160
rect 19475 5120 20076 5148
rect 19475 5117 19487 5120
rect 19429 5111 19487 5117
rect 20070 5108 20076 5120
rect 20128 5108 20134 5160
rect 15194 5080 15200 5092
rect 14844 5052 15200 5080
rect 14737 5043 14795 5049
rect 15194 5040 15200 5052
rect 15252 5080 15258 5092
rect 15838 5080 15844 5092
rect 15252 5052 15844 5080
rect 15252 5040 15258 5052
rect 15838 5040 15844 5052
rect 15896 5040 15902 5092
rect 16945 5083 17003 5089
rect 16945 5049 16957 5083
rect 16991 5080 17003 5083
rect 22020 5080 22048 5188
rect 22572 5157 22600 5188
rect 23106 5176 23112 5228
rect 23164 5176 23170 5228
rect 22373 5151 22431 5157
rect 22373 5117 22385 5151
rect 22419 5117 22431 5151
rect 22373 5111 22431 5117
rect 22557 5151 22615 5157
rect 22557 5117 22569 5151
rect 22603 5148 22615 5151
rect 22646 5148 22652 5160
rect 22603 5120 22652 5148
rect 22603 5117 22615 5120
rect 22557 5111 22615 5117
rect 16991 5052 22048 5080
rect 16991 5049 17003 5052
rect 16945 5043 17003 5049
rect 7006 4972 7012 5024
rect 7064 5012 7070 5024
rect 8113 5015 8171 5021
rect 8113 5012 8125 5015
rect 7064 4984 8125 5012
rect 7064 4972 7070 4984
rect 8113 4981 8125 4984
rect 8159 5012 8171 5015
rect 8478 5012 8484 5024
rect 8159 4984 8484 5012
rect 8159 4981 8171 4984
rect 8113 4975 8171 4981
rect 8478 4972 8484 4984
rect 8536 4972 8542 5024
rect 11974 4972 11980 5024
rect 12032 5012 12038 5024
rect 13357 5015 13415 5021
rect 13357 5012 13369 5015
rect 12032 4984 13369 5012
rect 12032 4972 12038 4984
rect 13357 4981 13369 4984
rect 13403 4981 13415 5015
rect 13357 4975 13415 4981
rect 13725 5015 13783 5021
rect 13725 4981 13737 5015
rect 13771 5012 13783 5015
rect 13814 5012 13820 5024
rect 13771 4984 13820 5012
rect 13771 4981 13783 4984
rect 13725 4975 13783 4981
rect 13814 4972 13820 4984
rect 13872 4972 13878 5024
rect 14461 5015 14519 5021
rect 14461 4981 14473 5015
rect 14507 5012 14519 5015
rect 14550 5012 14556 5024
rect 14507 4984 14556 5012
rect 14507 4981 14519 4984
rect 14461 4975 14519 4981
rect 14550 4972 14556 4984
rect 14608 4972 14614 5024
rect 20714 4972 20720 5024
rect 20772 5012 20778 5024
rect 21177 5015 21235 5021
rect 21177 5012 21189 5015
rect 20772 4984 21189 5012
rect 20772 4972 20778 4984
rect 21177 4981 21189 4984
rect 21223 4981 21235 5015
rect 22388 5012 22416 5111
rect 22646 5108 22652 5120
rect 22704 5108 22710 5160
rect 23385 5151 23443 5157
rect 23385 5148 23397 5151
rect 23124 5120 23397 5148
rect 23124 5092 23152 5120
rect 23385 5117 23397 5120
rect 23431 5117 23443 5151
rect 23385 5111 23443 5117
rect 23106 5040 23112 5092
rect 23164 5040 23170 5092
rect 24857 5015 24915 5021
rect 24857 5012 24869 5015
rect 22388 4984 24869 5012
rect 21177 4975 21235 4981
rect 24857 4981 24869 4984
rect 24903 5012 24915 5015
rect 24946 5012 24952 5024
rect 24903 4984 24952 5012
rect 24903 4981 24915 4984
rect 24857 4975 24915 4981
rect 24946 4972 24952 4984
rect 25004 4972 25010 5024
rect 1104 4922 25852 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 12214 4922
rect 12266 4870 12278 4922
rect 12330 4870 12342 4922
rect 12394 4870 12406 4922
rect 12458 4870 12470 4922
rect 12522 4870 20214 4922
rect 20266 4870 20278 4922
rect 20330 4870 20342 4922
rect 20394 4870 20406 4922
rect 20458 4870 20470 4922
rect 20522 4870 25852 4922
rect 1104 4848 25852 4870
rect 2501 4811 2559 4817
rect 2501 4777 2513 4811
rect 2547 4777 2559 4811
rect 2501 4771 2559 4777
rect 2685 4811 2743 4817
rect 2685 4777 2697 4811
rect 2731 4808 2743 4811
rect 3786 4808 3792 4820
rect 2731 4780 3792 4808
rect 2731 4777 2743 4780
rect 2685 4771 2743 4777
rect 2516 4740 2544 4771
rect 3786 4768 3792 4780
rect 3844 4768 3850 4820
rect 4111 4811 4169 4817
rect 4111 4777 4123 4811
rect 4157 4808 4169 4811
rect 4890 4808 4896 4820
rect 4157 4780 4896 4808
rect 4157 4777 4169 4780
rect 4111 4771 4169 4777
rect 4890 4768 4896 4780
rect 4948 4768 4954 4820
rect 5368 4780 7236 4808
rect 4985 4743 5043 4749
rect 2516 4712 4200 4740
rect 4172 4684 4200 4712
rect 4985 4709 4997 4743
rect 5031 4740 5043 4743
rect 5258 4740 5264 4752
rect 5031 4712 5264 4740
rect 5031 4709 5043 4712
rect 4985 4703 5043 4709
rect 5258 4700 5264 4712
rect 5316 4700 5322 4752
rect 2041 4675 2099 4681
rect 2041 4641 2053 4675
rect 2087 4672 2099 4675
rect 2498 4672 2504 4684
rect 2087 4644 2504 4672
rect 2087 4641 2099 4644
rect 2041 4635 2099 4641
rect 2498 4632 2504 4644
rect 2556 4632 2562 4684
rect 3050 4632 3056 4684
rect 3108 4672 3114 4684
rect 3237 4675 3295 4681
rect 3237 4672 3249 4675
rect 3108 4644 3249 4672
rect 3108 4632 3114 4644
rect 3237 4641 3249 4644
rect 3283 4641 3295 4675
rect 3237 4635 3295 4641
rect 3510 4632 3516 4684
rect 3568 4672 3574 4684
rect 3568 4644 4051 4672
rect 3568 4632 3574 4644
rect 1854 4564 1860 4616
rect 1912 4564 1918 4616
rect 3142 4604 3148 4616
rect 2332 4576 3148 4604
rect 2332 4545 2360 4576
rect 3142 4564 3148 4576
rect 3200 4564 3206 4616
rect 4023 4614 4051 4644
rect 4154 4632 4160 4684
rect 4212 4632 4218 4684
rect 4709 4675 4767 4681
rect 4709 4641 4721 4675
rect 4755 4672 4767 4675
rect 5368 4672 5396 4780
rect 5534 4700 5540 4752
rect 5592 4740 5598 4752
rect 5629 4743 5687 4749
rect 5629 4740 5641 4743
rect 5592 4712 5641 4740
rect 5592 4700 5598 4712
rect 5629 4709 5641 4712
rect 5675 4709 5687 4743
rect 5629 4703 5687 4709
rect 6549 4743 6607 4749
rect 6549 4709 6561 4743
rect 6595 4740 6607 4743
rect 7208 4740 7236 4780
rect 7650 4768 7656 4820
rect 7708 4808 7714 4820
rect 7837 4811 7895 4817
rect 7837 4808 7849 4811
rect 7708 4780 7849 4808
rect 7708 4768 7714 4780
rect 7837 4777 7849 4780
rect 7883 4777 7895 4811
rect 7837 4771 7895 4777
rect 7926 4768 7932 4820
rect 7984 4808 7990 4820
rect 8389 4811 8447 4817
rect 8389 4808 8401 4811
rect 7984 4780 8401 4808
rect 7984 4768 7990 4780
rect 8389 4777 8401 4780
rect 8435 4777 8447 4811
rect 8389 4771 8447 4777
rect 9122 4768 9128 4820
rect 9180 4808 9186 4820
rect 9217 4811 9275 4817
rect 9217 4808 9229 4811
rect 9180 4780 9229 4808
rect 9180 4768 9186 4780
rect 9217 4777 9229 4780
rect 9263 4777 9275 4811
rect 9217 4771 9275 4777
rect 11882 4768 11888 4820
rect 11940 4768 11946 4820
rect 12345 4811 12403 4817
rect 12345 4777 12357 4811
rect 12391 4808 12403 4811
rect 12618 4808 12624 4820
rect 12391 4780 12624 4808
rect 12391 4777 12403 4780
rect 12345 4771 12403 4777
rect 12618 4768 12624 4780
rect 12676 4768 12682 4820
rect 13814 4768 13820 4820
rect 13872 4808 13878 4820
rect 16669 4811 16727 4817
rect 13872 4780 16620 4808
rect 13872 4768 13878 4780
rect 6595 4712 7144 4740
rect 7208 4712 8432 4740
rect 6595 4709 6607 4712
rect 6549 4703 6607 4709
rect 7116 4681 7144 4712
rect 4755 4644 5396 4672
rect 6273 4675 6331 4681
rect 4755 4641 4767 4644
rect 4709 4635 4767 4641
rect 3329 4607 3387 4613
rect 3329 4573 3341 4607
rect 3375 4604 3387 4607
rect 4008 4608 4066 4614
rect 3375 4576 3740 4604
rect 3375 4573 3387 4576
rect 3329 4567 3387 4573
rect 2317 4539 2375 4545
rect 2317 4505 2329 4539
rect 2363 4505 2375 4539
rect 2317 4499 2375 4505
rect 2533 4539 2591 4545
rect 2533 4505 2545 4539
rect 2579 4536 2591 4539
rect 2579 4508 2774 4536
rect 2579 4505 2591 4508
rect 2533 4499 2591 4505
rect 2746 4468 2774 4508
rect 3712 4480 3740 4576
rect 4008 4574 4020 4608
rect 4054 4604 4066 4608
rect 4617 4607 4675 4613
rect 4617 4604 4629 4607
rect 4054 4576 4629 4604
rect 4054 4574 4066 4576
rect 4008 4568 4066 4574
rect 4617 4573 4629 4576
rect 4663 4604 4675 4607
rect 4798 4604 4804 4616
rect 4663 4576 4804 4604
rect 4663 4573 4675 4576
rect 4617 4567 4675 4573
rect 4798 4564 4804 4576
rect 4856 4564 4862 4616
rect 5276 4613 5304 4644
rect 6273 4641 6285 4675
rect 6319 4641 6331 4675
rect 6273 4635 6331 4641
rect 7101 4675 7159 4681
rect 7101 4641 7113 4675
rect 7147 4672 7159 4675
rect 8404 4672 8432 4712
rect 10502 4700 10508 4752
rect 10560 4700 10566 4752
rect 11146 4700 11152 4752
rect 11204 4740 11210 4752
rect 13832 4740 13860 4768
rect 11204 4712 13860 4740
rect 11204 4700 11210 4712
rect 16022 4700 16028 4752
rect 16080 4740 16086 4752
rect 16485 4743 16543 4749
rect 16485 4740 16497 4743
rect 16080 4712 16497 4740
rect 16080 4700 16086 4712
rect 16485 4709 16497 4712
rect 16531 4709 16543 4743
rect 16592 4740 16620 4780
rect 16669 4777 16681 4811
rect 16715 4808 16727 4811
rect 16942 4808 16948 4820
rect 16715 4780 16948 4808
rect 16715 4777 16727 4780
rect 16669 4771 16727 4777
rect 16942 4768 16948 4780
rect 17000 4768 17006 4820
rect 17126 4768 17132 4820
rect 17184 4808 17190 4820
rect 20898 4808 20904 4820
rect 17184 4780 20904 4808
rect 17184 4768 17190 4780
rect 19334 4740 19340 4752
rect 16592 4712 19340 4740
rect 16485 4703 16543 4709
rect 19334 4700 19340 4712
rect 19392 4700 19398 4752
rect 11974 4672 11980 4684
rect 7147 4644 8340 4672
rect 8404 4644 11980 4672
rect 7147 4641 7159 4644
rect 7101 4635 7159 4641
rect 5261 4607 5319 4613
rect 5261 4573 5273 4607
rect 5307 4573 5319 4607
rect 5261 4567 5319 4573
rect 5354 4607 5412 4613
rect 5354 4573 5366 4607
rect 5400 4573 5412 4607
rect 5354 4567 5412 4573
rect 6181 4607 6239 4613
rect 6181 4573 6193 4607
rect 6227 4573 6239 4607
rect 6181 4567 6239 4573
rect 4816 4536 4844 4564
rect 5369 4536 5397 4567
rect 4816 4508 5397 4536
rect 2961 4471 3019 4477
rect 2961 4468 2973 4471
rect 2746 4440 2973 4468
rect 2961 4437 2973 4440
rect 3007 4437 3019 4471
rect 2961 4431 3019 4437
rect 3694 4428 3700 4480
rect 3752 4468 3758 4480
rect 6196 4468 6224 4567
rect 6288 4536 6316 4635
rect 7006 4564 7012 4616
rect 7064 4564 7070 4616
rect 7190 4564 7196 4616
rect 7248 4604 7254 4616
rect 8312 4613 8340 4644
rect 11974 4632 11980 4644
rect 12032 4632 12038 4684
rect 13630 4672 13636 4684
rect 12360 4644 13636 4672
rect 7867 4607 7925 4613
rect 7867 4604 7879 4607
rect 7248 4576 7879 4604
rect 7248 4564 7254 4576
rect 7867 4573 7879 4576
rect 7913 4573 7925 4607
rect 7867 4567 7925 4573
rect 8021 4607 8079 4613
rect 8021 4573 8033 4607
rect 8067 4573 8079 4607
rect 8021 4567 8079 4573
rect 8297 4607 8355 4613
rect 8297 4573 8309 4607
rect 8343 4573 8355 4607
rect 8297 4567 8355 4573
rect 8036 4536 8064 4567
rect 8478 4564 8484 4616
rect 8536 4564 8542 4616
rect 9217 4607 9275 4613
rect 9217 4573 9229 4607
rect 9263 4604 9275 4607
rect 9306 4604 9312 4616
rect 9263 4576 9312 4604
rect 9263 4573 9275 4576
rect 9217 4567 9275 4573
rect 9306 4564 9312 4576
rect 9364 4564 9370 4616
rect 9401 4607 9459 4613
rect 9401 4573 9413 4607
rect 9447 4604 9459 4607
rect 9950 4604 9956 4616
rect 9447 4576 9956 4604
rect 9447 4573 9459 4576
rect 9401 4567 9459 4573
rect 9950 4564 9956 4576
rect 10008 4564 10014 4616
rect 11422 4604 11428 4616
rect 10612 4576 11428 4604
rect 10612 4536 10640 4576
rect 11422 4564 11428 4576
rect 11480 4564 11486 4616
rect 12066 4564 12072 4616
rect 12124 4564 12130 4616
rect 12360 4613 12388 4644
rect 12820 4613 12848 4644
rect 13630 4632 13636 4644
rect 13688 4632 13694 4684
rect 14185 4675 14243 4681
rect 14185 4641 14197 4675
rect 14231 4672 14243 4675
rect 14458 4672 14464 4684
rect 14231 4644 14464 4672
rect 14231 4641 14243 4644
rect 14185 4635 14243 4641
rect 14458 4632 14464 4644
rect 14516 4632 14522 4684
rect 18782 4632 18788 4684
rect 18840 4672 18846 4684
rect 19904 4681 19932 4780
rect 20898 4768 20904 4780
rect 20956 4808 20962 4820
rect 22189 4811 22247 4817
rect 20956 4780 22140 4808
rect 20956 4768 20962 4780
rect 22112 4740 22140 4780
rect 22189 4777 22201 4811
rect 22235 4808 22247 4811
rect 22370 4808 22376 4820
rect 22235 4780 22376 4808
rect 22235 4777 22247 4780
rect 22189 4771 22247 4777
rect 22370 4768 22376 4780
rect 22428 4768 22434 4820
rect 23106 4768 23112 4820
rect 23164 4768 23170 4820
rect 23382 4768 23388 4820
rect 23440 4768 23446 4820
rect 24854 4808 24860 4820
rect 23584 4780 24860 4808
rect 23584 4740 23612 4780
rect 24854 4768 24860 4780
rect 24912 4808 24918 4820
rect 24912 4780 24992 4808
rect 24912 4768 24918 4780
rect 22112 4712 23612 4740
rect 24489 4743 24547 4749
rect 24489 4709 24501 4743
rect 24535 4709 24547 4743
rect 24964 4740 24992 4780
rect 24964 4712 25084 4740
rect 24489 4703 24547 4709
rect 19889 4675 19947 4681
rect 18840 4644 19748 4672
rect 18840 4632 18846 4644
rect 12345 4607 12403 4613
rect 12345 4573 12357 4607
rect 12391 4573 12403 4607
rect 12345 4567 12403 4573
rect 12529 4607 12587 4613
rect 12529 4573 12541 4607
rect 12575 4573 12587 4607
rect 12529 4567 12587 4573
rect 12805 4607 12863 4613
rect 12805 4573 12817 4607
rect 12851 4573 12863 4607
rect 12805 4567 12863 4573
rect 12989 4607 13047 4613
rect 12989 4573 13001 4607
rect 13035 4573 13047 4607
rect 12989 4567 13047 4573
rect 6288 4508 10640 4536
rect 10689 4539 10747 4545
rect 10689 4505 10701 4539
rect 10735 4505 10747 4539
rect 12544 4536 12572 4567
rect 12618 4536 12624 4548
rect 12544 4508 12624 4536
rect 10689 4499 10747 4505
rect 7190 4468 7196 4480
rect 3752 4440 7196 4468
rect 3752 4428 3758 4440
rect 7190 4428 7196 4440
rect 7248 4428 7254 4480
rect 7377 4471 7435 4477
rect 7377 4437 7389 4471
rect 7423 4468 7435 4471
rect 7466 4468 7472 4480
rect 7423 4440 7472 4468
rect 7423 4437 7435 4440
rect 7377 4431 7435 4437
rect 7466 4428 7472 4440
rect 7524 4468 7530 4480
rect 8018 4468 8024 4480
rect 7524 4440 8024 4468
rect 7524 4428 7530 4440
rect 8018 4428 8024 4440
rect 8076 4428 8082 4480
rect 10704 4468 10732 4499
rect 12618 4496 12624 4508
rect 12676 4536 12682 4548
rect 13004 4536 13032 4567
rect 13722 4564 13728 4616
rect 13780 4564 13786 4616
rect 17678 4564 17684 4616
rect 17736 4564 17742 4616
rect 19720 4613 19748 4644
rect 19889 4641 19901 4675
rect 19935 4641 19947 4675
rect 19889 4635 19947 4641
rect 20714 4632 20720 4684
rect 20772 4632 20778 4684
rect 23750 4672 23756 4684
rect 22480 4644 23756 4672
rect 18693 4607 18751 4613
rect 18693 4573 18705 4607
rect 18739 4604 18751 4607
rect 19705 4607 19763 4613
rect 18739 4576 19380 4604
rect 18739 4573 18751 4576
rect 18693 4567 18751 4573
rect 13541 4539 13599 4545
rect 13541 4536 13553 4539
rect 12676 4508 13553 4536
rect 12676 4496 12682 4508
rect 13541 4505 13553 4508
rect 13587 4505 13599 4539
rect 13541 4499 13599 4505
rect 14366 4496 14372 4548
rect 14424 4536 14430 4548
rect 14461 4539 14519 4545
rect 14461 4536 14473 4539
rect 14424 4508 14473 4536
rect 14424 4496 14430 4508
rect 14461 4505 14473 4508
rect 14507 4505 14519 4539
rect 14461 4499 14519 4505
rect 14550 4496 14556 4548
rect 14608 4536 14614 4548
rect 14608 4508 14950 4536
rect 14608 4496 14614 4508
rect 16114 4496 16120 4548
rect 16172 4536 16178 4548
rect 16209 4539 16267 4545
rect 16209 4536 16221 4539
rect 16172 4508 16221 4536
rect 16172 4496 16178 4508
rect 16209 4505 16221 4508
rect 16255 4505 16267 4539
rect 16209 4499 16267 4505
rect 11514 4468 11520 4480
rect 10704 4440 11520 4468
rect 11514 4428 11520 4440
rect 11572 4428 11578 4480
rect 12897 4471 12955 4477
rect 12897 4437 12909 4471
rect 12943 4468 12955 4471
rect 12986 4468 12992 4480
rect 12943 4440 12992 4468
rect 12943 4437 12955 4440
rect 12897 4431 12955 4437
rect 12986 4428 12992 4440
rect 13044 4428 13050 4480
rect 15102 4428 15108 4480
rect 15160 4468 15166 4480
rect 15933 4471 15991 4477
rect 15933 4468 15945 4471
rect 15160 4440 15945 4468
rect 15160 4428 15166 4440
rect 15933 4437 15945 4440
rect 15979 4437 15991 4471
rect 15933 4431 15991 4437
rect 17494 4428 17500 4480
rect 17552 4428 17558 4480
rect 18506 4428 18512 4480
rect 18564 4428 18570 4480
rect 19352 4477 19380 4576
rect 19705 4573 19717 4607
rect 19751 4573 19763 4607
rect 19705 4567 19763 4573
rect 19794 4564 19800 4616
rect 19852 4604 19858 4616
rect 22480 4613 22508 4644
rect 23750 4632 23756 4644
rect 23808 4632 23814 4684
rect 23842 4632 23848 4684
rect 23900 4632 23906 4684
rect 24026 4632 24032 4684
rect 24084 4632 24090 4684
rect 20441 4607 20499 4613
rect 20441 4604 20453 4607
rect 19852 4576 20453 4604
rect 19852 4564 19858 4576
rect 20441 4573 20453 4576
rect 20487 4573 20499 4607
rect 20441 4567 20499 4573
rect 22465 4607 22523 4613
rect 22465 4573 22477 4607
rect 22511 4573 22523 4607
rect 22465 4567 22523 4573
rect 20990 4496 20996 4548
rect 21048 4536 21054 4548
rect 21048 4508 21206 4536
rect 21048 4496 21054 4508
rect 19337 4471 19395 4477
rect 19337 4437 19349 4471
rect 19383 4437 19395 4471
rect 19337 4431 19395 4437
rect 19797 4471 19855 4477
rect 19797 4437 19809 4471
rect 19843 4468 19855 4471
rect 19886 4468 19892 4480
rect 19843 4440 19892 4468
rect 19843 4437 19855 4440
rect 19797 4431 19855 4437
rect 19886 4428 19892 4440
rect 19944 4428 19950 4480
rect 20346 4428 20352 4480
rect 20404 4468 20410 4480
rect 22480 4468 22508 4567
rect 22554 4564 22560 4616
rect 22612 4604 22618 4616
rect 22649 4607 22707 4613
rect 22649 4604 22661 4607
rect 22612 4576 22661 4604
rect 22612 4564 22618 4576
rect 22649 4573 22661 4576
rect 22695 4573 22707 4607
rect 22649 4567 22707 4573
rect 22925 4607 22983 4613
rect 22925 4573 22937 4607
rect 22971 4604 22983 4607
rect 24504 4604 24532 4703
rect 24946 4632 24952 4684
rect 25004 4632 25010 4684
rect 25056 4681 25084 4712
rect 25041 4675 25099 4681
rect 25041 4641 25053 4675
rect 25087 4641 25099 4675
rect 25041 4635 25099 4641
rect 22971 4576 24532 4604
rect 22971 4573 22983 4576
rect 22925 4567 22983 4573
rect 20404 4440 22508 4468
rect 20404 4428 20410 4440
rect 22554 4428 22560 4480
rect 22612 4428 22618 4480
rect 23753 4471 23811 4477
rect 23753 4437 23765 4471
rect 23799 4468 23811 4471
rect 24762 4468 24768 4480
rect 23799 4440 24768 4468
rect 23799 4437 23811 4440
rect 23753 4431 23811 4437
rect 24762 4428 24768 4440
rect 24820 4468 24826 4480
rect 24857 4471 24915 4477
rect 24857 4468 24869 4471
rect 24820 4440 24869 4468
rect 24820 4428 24826 4440
rect 24857 4437 24869 4440
rect 24903 4437 24915 4471
rect 24857 4431 24915 4437
rect 1104 4378 25852 4400
rect 1104 4326 8214 4378
rect 8266 4326 8278 4378
rect 8330 4326 8342 4378
rect 8394 4326 8406 4378
rect 8458 4326 8470 4378
rect 8522 4326 16214 4378
rect 16266 4326 16278 4378
rect 16330 4326 16342 4378
rect 16394 4326 16406 4378
rect 16458 4326 16470 4378
rect 16522 4326 24214 4378
rect 24266 4326 24278 4378
rect 24330 4326 24342 4378
rect 24394 4326 24406 4378
rect 24458 4326 24470 4378
rect 24522 4326 25852 4378
rect 1104 4304 25852 4326
rect 4065 4267 4123 4273
rect 4065 4233 4077 4267
rect 4111 4264 4123 4267
rect 4154 4264 4160 4276
rect 4111 4236 4160 4264
rect 4111 4233 4123 4236
rect 4065 4227 4123 4233
rect 4154 4224 4160 4236
rect 4212 4224 4218 4276
rect 4249 4267 4307 4273
rect 4249 4233 4261 4267
rect 4295 4264 4307 4267
rect 4614 4264 4620 4276
rect 4295 4236 4620 4264
rect 4295 4233 4307 4236
rect 4249 4227 4307 4233
rect 4614 4224 4620 4236
rect 4672 4224 4678 4276
rect 6825 4267 6883 4273
rect 6825 4233 6837 4267
rect 6871 4264 6883 4267
rect 7190 4264 7196 4276
rect 6871 4236 7196 4264
rect 6871 4233 6883 4236
rect 6825 4227 6883 4233
rect 7190 4224 7196 4236
rect 7248 4224 7254 4276
rect 10137 4267 10195 4273
rect 7760 4236 8340 4264
rect 2958 4156 2964 4208
rect 3016 4156 3022 4208
rect 1486 4088 1492 4140
rect 1544 4128 1550 4140
rect 1673 4131 1731 4137
rect 1673 4128 1685 4131
rect 1544 4100 1685 4128
rect 1544 4088 1550 4100
rect 1673 4097 1685 4100
rect 1719 4097 1731 4131
rect 3694 4128 3700 4140
rect 1673 4091 1731 4097
rect 3436 4100 3700 4128
rect 1946 4020 1952 4072
rect 2004 4020 2010 4072
rect 3436 4069 3464 4100
rect 3694 4088 3700 4100
rect 3752 4088 3758 4140
rect 4172 4128 4200 4224
rect 4525 4131 4583 4137
rect 4525 4128 4537 4131
rect 4172 4100 4537 4128
rect 4525 4097 4537 4100
rect 4571 4097 4583 4131
rect 4798 4128 4804 4140
rect 4759 4100 4804 4128
rect 4525 4091 4583 4097
rect 4798 4088 4804 4100
rect 4856 4088 4862 4140
rect 4893 4131 4951 4137
rect 4893 4097 4905 4131
rect 4939 4128 4951 4131
rect 4982 4128 4988 4140
rect 4939 4100 4988 4128
rect 4939 4097 4951 4100
rect 4893 4091 4951 4097
rect 4982 4088 4988 4100
rect 5040 4088 5046 4140
rect 7466 4088 7472 4140
rect 7524 4088 7530 4140
rect 7760 4137 7788 4236
rect 8018 4156 8024 4208
rect 8076 4156 8082 4208
rect 7561 4131 7619 4137
rect 7561 4097 7573 4131
rect 7607 4097 7619 4131
rect 7561 4091 7619 4097
rect 7745 4131 7803 4137
rect 7745 4097 7757 4131
rect 7791 4097 7803 4131
rect 7745 4091 7803 4097
rect 3421 4063 3479 4069
rect 3421 4029 3433 4063
rect 3467 4029 3479 4063
rect 3421 4023 3479 4029
rect 6638 4020 6644 4072
rect 6696 4060 6702 4072
rect 6917 4063 6975 4069
rect 6917 4060 6929 4063
rect 6696 4032 6929 4060
rect 6696 4020 6702 4032
rect 6917 4029 6929 4032
rect 6963 4029 6975 4063
rect 6917 4023 6975 4029
rect 7098 4020 7104 4072
rect 7156 4020 7162 4072
rect 7576 4060 7604 4091
rect 8110 4088 8116 4140
rect 8168 4128 8174 4140
rect 8312 4137 8340 4236
rect 10137 4233 10149 4267
rect 10183 4264 10195 4267
rect 10502 4264 10508 4276
rect 10183 4236 10508 4264
rect 10183 4233 10195 4236
rect 10137 4227 10195 4233
rect 10502 4224 10508 4236
rect 10560 4224 10566 4276
rect 10962 4224 10968 4276
rect 11020 4264 11026 4276
rect 14458 4264 14464 4276
rect 11020 4236 14464 4264
rect 11020 4224 11026 4236
rect 10612 4168 10824 4196
rect 10612 4140 10640 4168
rect 8205 4131 8263 4137
rect 8205 4128 8217 4131
rect 8168 4100 8217 4128
rect 8168 4088 8174 4100
rect 8205 4097 8217 4100
rect 8251 4097 8263 4131
rect 8205 4091 8263 4097
rect 8297 4131 8355 4137
rect 8297 4097 8309 4131
rect 8343 4128 8355 4131
rect 8570 4128 8576 4140
rect 8343 4100 8576 4128
rect 8343 4097 8355 4100
rect 8297 4091 8355 4097
rect 8570 4088 8576 4100
rect 8628 4088 8634 4140
rect 8662 4088 8668 4140
rect 8720 4128 8726 4140
rect 9122 4128 9128 4140
rect 8720 4100 9128 4128
rect 8720 4088 8726 4100
rect 9122 4088 9128 4100
rect 9180 4088 9186 4140
rect 9953 4131 10011 4137
rect 9953 4128 9965 4131
rect 9324 4100 9965 4128
rect 8128 4060 8156 4088
rect 7576 4032 8156 4060
rect 9214 4020 9220 4072
rect 9272 4020 9278 4072
rect 3050 3952 3056 4004
rect 3108 3992 3114 4004
rect 3108 3964 3556 3992
rect 3108 3952 3114 3964
rect 3528 3924 3556 3964
rect 6270 3952 6276 4004
rect 6328 3992 6334 4004
rect 6328 3964 7604 3992
rect 6328 3952 6334 3964
rect 7576 3936 7604 3964
rect 8294 3952 8300 4004
rect 8352 3992 8358 4004
rect 8754 3992 8760 4004
rect 8352 3964 8760 3992
rect 8352 3952 8358 3964
rect 8754 3952 8760 3964
rect 8812 3992 8818 4004
rect 9324 3992 9352 4100
rect 9953 4097 9965 4100
rect 9999 4097 10011 4131
rect 9953 4091 10011 4097
rect 10229 4131 10287 4137
rect 10229 4097 10241 4131
rect 10275 4097 10287 4131
rect 10229 4091 10287 4097
rect 10505 4131 10563 4137
rect 10505 4097 10517 4131
rect 10551 4128 10563 4131
rect 10594 4128 10600 4140
rect 10551 4100 10600 4128
rect 10551 4097 10563 4100
rect 10505 4091 10563 4097
rect 9493 4063 9551 4069
rect 9493 4029 9505 4063
rect 9539 4060 9551 4063
rect 10244 4060 10272 4091
rect 10594 4088 10600 4100
rect 10652 4088 10658 4140
rect 10689 4131 10747 4137
rect 10689 4097 10701 4131
rect 10735 4097 10747 4131
rect 10796 4128 10824 4168
rect 10965 4131 11023 4137
rect 10965 4128 10977 4131
rect 10796 4100 10977 4128
rect 10689 4091 10747 4097
rect 10965 4097 10977 4100
rect 11011 4097 11023 4131
rect 10965 4091 11023 4097
rect 9539 4032 10272 4060
rect 10704 4060 10732 4091
rect 11146 4088 11152 4140
rect 11204 4088 11210 4140
rect 11716 4137 11744 4236
rect 14458 4224 14464 4236
rect 14516 4224 14522 4276
rect 17497 4267 17555 4273
rect 17497 4233 17509 4267
rect 17543 4264 17555 4267
rect 17586 4264 17592 4276
rect 17543 4236 17592 4264
rect 17543 4233 17555 4236
rect 17497 4227 17555 4233
rect 17586 4224 17592 4236
rect 17644 4224 17650 4276
rect 17678 4224 17684 4276
rect 17736 4264 17742 4276
rect 17865 4267 17923 4273
rect 17865 4264 17877 4267
rect 17736 4236 17877 4264
rect 17736 4224 17742 4236
rect 17865 4233 17877 4236
rect 17911 4233 17923 4267
rect 17865 4227 17923 4233
rect 19334 4224 19340 4276
rect 19392 4264 19398 4276
rect 20622 4264 20628 4276
rect 19392 4236 20628 4264
rect 19392 4224 19398 4236
rect 12986 4156 12992 4208
rect 13044 4156 13050 4208
rect 16482 4196 16488 4208
rect 16146 4168 16488 4196
rect 16482 4156 16488 4168
rect 16540 4156 16546 4208
rect 18417 4199 18475 4205
rect 18417 4165 18429 4199
rect 18463 4196 18475 4199
rect 18506 4196 18512 4208
rect 18463 4168 18512 4196
rect 18463 4165 18475 4168
rect 18417 4159 18475 4165
rect 18506 4156 18512 4168
rect 18564 4156 18570 4208
rect 11701 4131 11759 4137
rect 11701 4097 11713 4131
rect 11747 4097 11759 4131
rect 11701 4091 11759 4097
rect 14182 4088 14188 4140
rect 14240 4088 14246 4140
rect 14458 4088 14464 4140
rect 14516 4128 14522 4140
rect 20180 4137 20208 4236
rect 20622 4224 20628 4236
rect 20680 4224 20686 4276
rect 24762 4224 24768 4276
rect 24820 4224 24826 4276
rect 22554 4156 22560 4208
rect 22612 4196 22618 4208
rect 22612 4168 23782 4196
rect 22612 4156 22618 4168
rect 14645 4131 14703 4137
rect 14645 4128 14657 4131
rect 14516 4100 14657 4128
rect 14516 4088 14522 4100
rect 14645 4097 14657 4100
rect 14691 4097 14703 4131
rect 20165 4131 20223 4137
rect 14645 4091 14703 4097
rect 11164 4060 11192 4088
rect 10704 4032 11192 4060
rect 9539 4029 9551 4032
rect 9493 4023 9551 4029
rect 11974 4020 11980 4072
rect 12032 4020 12038 4072
rect 14921 4063 14979 4069
rect 14921 4029 14933 4063
rect 14967 4060 14979 4063
rect 16114 4060 16120 4072
rect 14967 4032 16120 4060
rect 14967 4029 14979 4032
rect 14921 4023 14979 4029
rect 16114 4020 16120 4032
rect 16172 4060 16178 4072
rect 16172 4032 16574 4060
rect 16172 4020 16178 4032
rect 11330 3992 11336 4004
rect 8812 3964 9352 3992
rect 9416 3964 11336 3992
rect 8812 3952 8818 3964
rect 4065 3927 4123 3933
rect 4065 3924 4077 3927
rect 3528 3896 4077 3924
rect 4065 3893 4077 3896
rect 4111 3893 4123 3927
rect 4065 3887 4123 3893
rect 4798 3884 4804 3936
rect 4856 3924 4862 3936
rect 6457 3927 6515 3933
rect 6457 3924 6469 3927
rect 4856 3896 6469 3924
rect 4856 3884 4862 3896
rect 6457 3893 6469 3896
rect 6503 3893 6515 3927
rect 6457 3887 6515 3893
rect 7466 3884 7472 3936
rect 7524 3884 7530 3936
rect 7558 3884 7564 3936
rect 7616 3924 7622 3936
rect 8021 3927 8079 3933
rect 8021 3924 8033 3927
rect 7616 3896 8033 3924
rect 7616 3884 7622 3896
rect 8021 3893 8033 3896
rect 8067 3893 8079 3927
rect 8021 3887 8079 3893
rect 9122 3884 9128 3936
rect 9180 3924 9186 3936
rect 9416 3924 9444 3964
rect 11330 3952 11336 3964
rect 11388 3952 11394 4004
rect 14366 3952 14372 4004
rect 14424 3952 14430 4004
rect 16022 3952 16028 4004
rect 16080 3992 16086 4004
rect 16393 3995 16451 4001
rect 16393 3992 16405 3995
rect 16080 3964 16405 3992
rect 16080 3952 16086 3964
rect 16393 3961 16405 3964
rect 16439 3961 16451 3995
rect 16393 3955 16451 3961
rect 9180 3896 9444 3924
rect 9180 3884 9186 3896
rect 9766 3884 9772 3936
rect 9824 3884 9830 3936
rect 10594 3884 10600 3936
rect 10652 3924 10658 3936
rect 10689 3927 10747 3933
rect 10689 3924 10701 3927
rect 10652 3896 10701 3924
rect 10652 3884 10658 3896
rect 10689 3893 10701 3896
rect 10735 3893 10747 3927
rect 10689 3887 10747 3893
rect 11146 3884 11152 3936
rect 11204 3884 11210 3936
rect 11422 3884 11428 3936
rect 11480 3924 11486 3936
rect 12986 3924 12992 3936
rect 11480 3896 12992 3924
rect 11480 3884 11486 3896
rect 12986 3884 12992 3896
rect 13044 3924 13050 3936
rect 13449 3927 13507 3933
rect 13449 3924 13461 3927
rect 13044 3896 13461 3924
rect 13044 3884 13050 3896
rect 13449 3893 13461 3896
rect 13495 3893 13507 3927
rect 16546 3924 16574 4032
rect 17126 4020 17132 4072
rect 17184 4060 17190 4072
rect 17221 4063 17279 4069
rect 17221 4060 17233 4063
rect 17184 4032 17233 4060
rect 17184 4020 17190 4032
rect 17221 4029 17233 4032
rect 17267 4029 17279 4063
rect 17221 4023 17279 4029
rect 17405 4063 17463 4069
rect 17405 4029 17417 4063
rect 17451 4060 17463 4063
rect 17586 4060 17592 4072
rect 17451 4032 17592 4060
rect 17451 4029 17463 4032
rect 17405 4023 17463 4029
rect 17586 4020 17592 4032
rect 17644 4020 17650 4072
rect 18141 4063 18199 4069
rect 18141 4029 18153 4063
rect 18187 4029 18199 4063
rect 19536 4060 19564 4114
rect 20165 4097 20177 4131
rect 20211 4097 20223 4131
rect 20165 4091 20223 4097
rect 20346 4088 20352 4140
rect 20404 4088 20410 4140
rect 20806 4088 20812 4140
rect 20864 4088 20870 4140
rect 20993 4131 21051 4137
rect 20993 4128 21005 4131
rect 20916 4100 21005 4128
rect 20257 4063 20315 4069
rect 20257 4060 20269 4063
rect 19536 4032 20269 4060
rect 18141 4023 18199 4029
rect 20257 4029 20269 4032
rect 20303 4029 20315 4063
rect 20257 4023 20315 4029
rect 16666 3952 16672 4004
rect 16724 3992 16730 4004
rect 18156 3992 18184 4023
rect 16724 3964 18184 3992
rect 16724 3952 16730 3964
rect 18046 3924 18052 3936
rect 16546 3896 18052 3924
rect 13449 3887 13507 3893
rect 18046 3884 18052 3896
rect 18104 3884 18110 3936
rect 18156 3924 18184 3964
rect 19610 3952 19616 4004
rect 19668 3992 19674 4004
rect 20916 3992 20944 4100
rect 20993 4097 21005 4100
rect 21039 4097 21051 4131
rect 20993 4091 21051 4097
rect 23014 4088 23020 4140
rect 23072 4088 23078 4140
rect 23290 4020 23296 4072
rect 23348 4020 23354 4072
rect 19668 3964 20944 3992
rect 19668 3952 19674 3964
rect 20990 3952 20996 4004
rect 21048 3952 21054 4004
rect 19794 3924 19800 3936
rect 18156 3896 19800 3924
rect 19794 3884 19800 3896
rect 19852 3884 19858 3936
rect 19886 3884 19892 3936
rect 19944 3884 19950 3936
rect 1104 3834 25852 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 12214 3834
rect 12266 3782 12278 3834
rect 12330 3782 12342 3834
rect 12394 3782 12406 3834
rect 12458 3782 12470 3834
rect 12522 3782 20214 3834
rect 20266 3782 20278 3834
rect 20330 3782 20342 3834
rect 20394 3782 20406 3834
rect 20458 3782 20470 3834
rect 20522 3782 25852 3834
rect 1104 3760 25852 3782
rect 1946 3680 1952 3732
rect 2004 3720 2010 3732
rect 2225 3723 2283 3729
rect 2225 3720 2237 3723
rect 2004 3692 2237 3720
rect 2004 3680 2010 3692
rect 2225 3689 2237 3692
rect 2271 3689 2283 3723
rect 2225 3683 2283 3689
rect 2777 3723 2835 3729
rect 2777 3689 2789 3723
rect 2823 3720 2835 3723
rect 2958 3720 2964 3732
rect 2823 3692 2964 3720
rect 2823 3689 2835 3692
rect 2777 3683 2835 3689
rect 2958 3680 2964 3692
rect 3016 3680 3022 3732
rect 6638 3680 6644 3732
rect 6696 3680 6702 3732
rect 7374 3680 7380 3732
rect 7432 3680 7438 3732
rect 8846 3720 8852 3732
rect 8496 3692 8852 3720
rect 6178 3612 6184 3664
rect 6236 3652 6242 3664
rect 7466 3652 7472 3664
rect 6236 3624 7472 3652
rect 6236 3612 6242 3624
rect 7466 3612 7472 3624
rect 7524 3652 7530 3664
rect 7524 3624 7880 3652
rect 7524 3612 7530 3624
rect 4798 3584 4804 3596
rect 2424 3556 4804 3584
rect 2424 3525 2452 3556
rect 4798 3544 4804 3556
rect 4856 3544 4862 3596
rect 5905 3587 5963 3593
rect 5905 3553 5917 3587
rect 5951 3584 5963 3587
rect 7009 3587 7067 3593
rect 7009 3584 7021 3587
rect 5951 3556 7021 3584
rect 5951 3553 5963 3556
rect 5905 3547 5963 3553
rect 7009 3553 7021 3556
rect 7055 3553 7067 3587
rect 7009 3547 7067 3553
rect 2409 3519 2467 3525
rect 2409 3485 2421 3519
rect 2455 3485 2467 3519
rect 2409 3479 2467 3485
rect 2777 3519 2835 3525
rect 2777 3485 2789 3519
rect 2823 3516 2835 3519
rect 2866 3516 2872 3528
rect 2823 3488 2872 3516
rect 2823 3485 2835 3488
rect 2777 3479 2835 3485
rect 2866 3476 2872 3488
rect 2924 3476 2930 3528
rect 2961 3519 3019 3525
rect 2961 3485 2973 3519
rect 3007 3516 3019 3519
rect 4433 3519 4491 3525
rect 4433 3516 4445 3519
rect 3007 3488 4445 3516
rect 3007 3485 3019 3488
rect 2961 3479 3019 3485
rect 4433 3485 4445 3488
rect 4479 3485 4491 3519
rect 4433 3479 4491 3485
rect 4617 3519 4675 3525
rect 4617 3485 4629 3519
rect 4663 3485 4675 3519
rect 4617 3479 4675 3485
rect 2498 3408 2504 3460
rect 2556 3448 2562 3460
rect 2976 3448 3004 3479
rect 4632 3448 4660 3479
rect 6178 3476 6184 3528
rect 6236 3476 6242 3528
rect 6270 3476 6276 3528
rect 6328 3476 6334 3528
rect 6891 3519 6949 3525
rect 6891 3485 6903 3519
rect 6937 3516 6949 3519
rect 6937 3512 6960 3516
rect 6937 3485 7052 3512
rect 6891 3484 7052 3485
rect 6891 3479 6949 3484
rect 2556 3420 3004 3448
rect 4448 3420 4660 3448
rect 7024 3448 7052 3484
rect 7558 3476 7564 3528
rect 7616 3476 7622 3528
rect 7742 3476 7748 3528
rect 7800 3476 7806 3528
rect 7852 3525 7880 3624
rect 8496 3584 8524 3692
rect 8846 3680 8852 3692
rect 8904 3720 8910 3732
rect 10502 3720 10508 3732
rect 8904 3692 10508 3720
rect 8904 3680 8910 3692
rect 10502 3680 10508 3692
rect 10560 3680 10566 3732
rect 10965 3723 11023 3729
rect 10965 3689 10977 3723
rect 11011 3720 11023 3723
rect 11330 3720 11336 3732
rect 11011 3692 11336 3720
rect 11011 3689 11023 3692
rect 10965 3683 11023 3689
rect 11330 3680 11336 3692
rect 11388 3680 11394 3732
rect 11974 3680 11980 3732
rect 12032 3720 12038 3732
rect 12253 3723 12311 3729
rect 12253 3720 12265 3723
rect 12032 3692 12265 3720
rect 12032 3680 12038 3692
rect 12253 3689 12265 3692
rect 12299 3689 12311 3723
rect 12253 3683 12311 3689
rect 16482 3680 16488 3732
rect 16540 3680 16546 3732
rect 17586 3680 17592 3732
rect 17644 3720 17650 3732
rect 18969 3723 19027 3729
rect 18969 3720 18981 3723
rect 17644 3692 18981 3720
rect 17644 3680 17650 3692
rect 18969 3689 18981 3692
rect 19015 3689 19027 3723
rect 18969 3683 19027 3689
rect 20622 3680 20628 3732
rect 20680 3720 20686 3732
rect 23569 3723 23627 3729
rect 20680 3692 23152 3720
rect 20680 3680 20686 3692
rect 12713 3655 12771 3661
rect 12713 3621 12725 3655
rect 12759 3621 12771 3655
rect 12713 3615 12771 3621
rect 8404 3556 8524 3584
rect 7837 3519 7895 3525
rect 7837 3485 7849 3519
rect 7883 3485 7895 3519
rect 7837 3479 7895 3485
rect 8294 3476 8300 3528
rect 8352 3476 8358 3528
rect 8404 3525 8432 3556
rect 9030 3544 9036 3596
rect 9088 3584 9094 3596
rect 9217 3587 9275 3593
rect 9217 3584 9229 3587
rect 9088 3556 9229 3584
rect 9088 3544 9094 3556
rect 9217 3553 9229 3556
rect 9263 3584 9275 3587
rect 9858 3584 9864 3596
rect 9263 3556 9864 3584
rect 9263 3553 9275 3556
rect 9217 3547 9275 3553
rect 9858 3544 9864 3556
rect 9916 3584 9922 3596
rect 10962 3584 10968 3596
rect 9916 3556 10968 3584
rect 9916 3544 9922 3556
rect 10962 3544 10968 3556
rect 11020 3544 11026 3596
rect 8389 3519 8447 3525
rect 8389 3485 8401 3519
rect 8435 3485 8447 3519
rect 8389 3479 8447 3485
rect 8481 3519 8539 3525
rect 8481 3485 8493 3519
rect 8527 3485 8539 3519
rect 8481 3479 8539 3485
rect 7760 3448 7788 3476
rect 7024 3420 7788 3448
rect 8496 3448 8524 3479
rect 10594 3476 10600 3528
rect 10652 3476 10658 3528
rect 12437 3519 12495 3525
rect 12437 3485 12449 3519
rect 12483 3516 12495 3519
rect 12728 3516 12756 3615
rect 13078 3612 13084 3664
rect 13136 3652 13142 3664
rect 16666 3652 16672 3664
rect 13136 3624 14688 3652
rect 13136 3612 13142 3624
rect 13262 3544 13268 3596
rect 13320 3544 13326 3596
rect 12483 3488 12756 3516
rect 12483 3485 12495 3488
rect 12437 3479 12495 3485
rect 12986 3476 12992 3528
rect 13044 3516 13050 3528
rect 13081 3519 13139 3525
rect 13081 3516 13093 3519
rect 13044 3488 13093 3516
rect 13044 3476 13050 3488
rect 13081 3485 13093 3488
rect 13127 3485 13139 3519
rect 13081 3479 13139 3485
rect 9214 3448 9220 3460
rect 8496 3420 9220 3448
rect 2556 3408 2562 3420
rect 2866 3340 2872 3392
rect 2924 3380 2930 3392
rect 3602 3380 3608 3392
rect 2924 3352 3608 3380
rect 2924 3340 2930 3352
rect 3602 3340 3608 3352
rect 3660 3380 3666 3392
rect 4448 3380 4476 3420
rect 9214 3408 9220 3420
rect 9272 3408 9278 3460
rect 9493 3451 9551 3457
rect 9493 3417 9505 3451
rect 9539 3448 9551 3451
rect 9766 3448 9772 3460
rect 9539 3420 9772 3448
rect 9539 3417 9551 3420
rect 9493 3411 9551 3417
rect 9766 3408 9772 3420
rect 9824 3408 9830 3460
rect 12066 3408 12072 3460
rect 12124 3448 12130 3460
rect 13280 3448 13308 3544
rect 14185 3519 14243 3525
rect 14185 3485 14197 3519
rect 14231 3516 14243 3519
rect 14550 3516 14556 3528
rect 14231 3488 14556 3516
rect 14231 3485 14243 3488
rect 14185 3479 14243 3485
rect 14550 3476 14556 3488
rect 14608 3476 14614 3528
rect 14660 3516 14688 3624
rect 16546 3624 16672 3652
rect 15930 3544 15936 3596
rect 15988 3584 15994 3596
rect 16546 3584 16574 3624
rect 16666 3612 16672 3624
rect 16724 3612 16730 3664
rect 20717 3655 20775 3661
rect 20717 3621 20729 3655
rect 20763 3652 20775 3655
rect 21082 3652 21088 3664
rect 20763 3624 21088 3652
rect 20763 3621 20775 3624
rect 20717 3615 20775 3621
rect 21082 3612 21088 3624
rect 21140 3612 21146 3664
rect 17221 3587 17279 3593
rect 17221 3584 17233 3587
rect 15988 3556 17233 3584
rect 15988 3544 15994 3556
rect 17221 3553 17233 3556
rect 17267 3553 17279 3587
rect 17221 3547 17279 3553
rect 17494 3544 17500 3596
rect 17552 3544 17558 3596
rect 18046 3544 18052 3596
rect 18104 3584 18110 3596
rect 20993 3587 21051 3593
rect 20993 3584 21005 3587
rect 18104 3556 21005 3584
rect 18104 3544 18110 3556
rect 20993 3553 21005 3556
rect 21039 3553 21051 3587
rect 20993 3547 21051 3553
rect 22741 3587 22799 3593
rect 22741 3553 22753 3587
rect 22787 3584 22799 3587
rect 23014 3584 23020 3596
rect 22787 3556 23020 3584
rect 22787 3553 22799 3556
rect 22741 3547 22799 3553
rect 23014 3544 23020 3556
rect 23072 3544 23078 3596
rect 16485 3519 16543 3525
rect 16485 3516 16497 3519
rect 14660 3488 16497 3516
rect 16485 3485 16497 3488
rect 16531 3516 16543 3519
rect 16531 3488 16620 3516
rect 16531 3485 16543 3488
rect 16485 3479 16543 3485
rect 12124 3420 13308 3448
rect 12124 3408 12130 3420
rect 3660 3352 4476 3380
rect 4525 3383 4583 3389
rect 3660 3340 3666 3352
rect 4525 3349 4537 3383
rect 4571 3380 4583 3383
rect 4614 3380 4620 3392
rect 4571 3352 4620 3380
rect 4571 3349 4583 3352
rect 4525 3343 4583 3349
rect 4614 3340 4620 3352
rect 4672 3340 4678 3392
rect 8665 3383 8723 3389
rect 8665 3349 8677 3383
rect 8711 3380 8723 3383
rect 9306 3380 9312 3392
rect 8711 3352 9312 3380
rect 8711 3349 8723 3352
rect 8665 3343 8723 3349
rect 9306 3340 9312 3352
rect 9364 3340 9370 3392
rect 13173 3383 13231 3389
rect 13173 3349 13185 3383
rect 13219 3380 13231 3383
rect 14182 3380 14188 3392
rect 13219 3352 14188 3380
rect 13219 3349 13231 3352
rect 13173 3343 13231 3349
rect 14182 3340 14188 3352
rect 14240 3340 14246 3392
rect 14369 3383 14427 3389
rect 14369 3349 14381 3383
rect 14415 3380 14427 3383
rect 15010 3380 15016 3392
rect 14415 3352 15016 3380
rect 14415 3349 14427 3352
rect 14369 3343 14427 3349
rect 15010 3340 15016 3352
rect 15068 3340 15074 3392
rect 16592 3380 16620 3488
rect 16666 3476 16672 3528
rect 16724 3476 16730 3528
rect 19334 3476 19340 3528
rect 19392 3476 19398 3528
rect 19521 3519 19579 3525
rect 19521 3485 19533 3519
rect 19567 3516 19579 3519
rect 20070 3516 20076 3528
rect 19567 3488 20076 3516
rect 19567 3485 19579 3488
rect 19521 3479 19579 3485
rect 20070 3476 20076 3488
rect 20128 3476 20134 3528
rect 20533 3519 20591 3525
rect 20533 3485 20545 3519
rect 20579 3485 20591 3519
rect 20533 3479 20591 3485
rect 20717 3519 20775 3525
rect 20717 3485 20729 3519
rect 20763 3485 20775 3519
rect 23124 3516 23152 3692
rect 23569 3689 23581 3723
rect 23615 3720 23627 3723
rect 23658 3720 23664 3732
rect 23615 3692 23664 3720
rect 23615 3689 23627 3692
rect 23569 3683 23627 3689
rect 23658 3680 23664 3692
rect 23716 3680 23722 3732
rect 23566 3516 23572 3528
rect 23124 3488 23572 3516
rect 20717 3479 20775 3485
rect 19429 3451 19487 3457
rect 19429 3448 19441 3451
rect 18722 3420 19441 3448
rect 19429 3417 19441 3420
rect 19475 3417 19487 3451
rect 19429 3411 19487 3417
rect 19702 3408 19708 3460
rect 19760 3448 19766 3460
rect 20548 3448 20576 3479
rect 20622 3448 20628 3460
rect 19760 3420 20628 3448
rect 19760 3408 19766 3420
rect 20622 3408 20628 3420
rect 20680 3408 20686 3460
rect 20732 3380 20760 3479
rect 23566 3476 23572 3488
rect 23624 3476 23630 3528
rect 23750 3476 23756 3528
rect 23808 3476 23814 3528
rect 22002 3408 22008 3460
rect 22060 3408 22066 3460
rect 22465 3451 22523 3457
rect 22465 3417 22477 3451
rect 22511 3417 22523 3451
rect 22465 3411 22523 3417
rect 21450 3380 21456 3392
rect 16592 3352 21456 3380
rect 21450 3340 21456 3352
rect 21508 3340 21514 3392
rect 21542 3340 21548 3392
rect 21600 3380 21606 3392
rect 22480 3380 22508 3411
rect 21600 3352 22508 3380
rect 21600 3340 21606 3352
rect 1104 3290 25852 3312
rect 1104 3238 8214 3290
rect 8266 3238 8278 3290
rect 8330 3238 8342 3290
rect 8394 3238 8406 3290
rect 8458 3238 8470 3290
rect 8522 3238 16214 3290
rect 16266 3238 16278 3290
rect 16330 3238 16342 3290
rect 16394 3238 16406 3290
rect 16458 3238 16470 3290
rect 16522 3238 24214 3290
rect 24266 3238 24278 3290
rect 24330 3238 24342 3290
rect 24394 3238 24406 3290
rect 24458 3238 24470 3290
rect 24522 3238 25852 3290
rect 1104 3216 25852 3238
rect 3881 3179 3939 3185
rect 3881 3145 3893 3179
rect 3927 3176 3939 3179
rect 4706 3176 4712 3188
rect 3927 3148 4712 3176
rect 3927 3145 3939 3148
rect 3881 3139 3939 3145
rect 4706 3136 4712 3148
rect 4764 3136 4770 3188
rect 5166 3136 5172 3188
rect 5224 3176 5230 3188
rect 5261 3179 5319 3185
rect 5261 3176 5273 3179
rect 5224 3148 5273 3176
rect 5224 3136 5230 3148
rect 5261 3145 5273 3148
rect 5307 3145 5319 3179
rect 7653 3179 7711 3185
rect 7653 3176 7665 3179
rect 5261 3139 5319 3145
rect 5736 3148 7665 3176
rect 4249 3111 4307 3117
rect 4249 3077 4261 3111
rect 4295 3108 4307 3111
rect 4893 3111 4951 3117
rect 4893 3108 4905 3111
rect 4295 3080 4905 3108
rect 4295 3077 4307 3080
rect 4249 3071 4307 3077
rect 4893 3077 4905 3080
rect 4939 3108 4951 3111
rect 5537 3111 5595 3117
rect 5537 3108 5549 3111
rect 4939 3080 5549 3108
rect 4939 3077 4951 3080
rect 4893 3071 4951 3077
rect 5537 3077 5549 3080
rect 5583 3077 5595 3111
rect 5537 3071 5595 3077
rect 2498 3000 2504 3052
rect 2556 3040 2562 3052
rect 3421 3043 3479 3049
rect 3421 3040 3433 3043
rect 2556 3012 3433 3040
rect 2556 3000 2562 3012
rect 3421 3009 3433 3012
rect 3467 3009 3479 3043
rect 3421 3003 3479 3009
rect 3602 3000 3608 3052
rect 3660 3000 3666 3052
rect 4065 3043 4123 3049
rect 4065 3009 4077 3043
rect 4111 3009 4123 3043
rect 4065 3003 4123 3009
rect 4341 3043 4399 3049
rect 4341 3009 4353 3043
rect 4387 3040 4399 3043
rect 4387 3012 5028 3040
rect 4387 3009 4399 3012
rect 4341 3003 4399 3009
rect 4080 2972 4108 3003
rect 5000 2984 5028 3012
rect 4617 2975 4675 2981
rect 4617 2972 4629 2975
rect 4080 2944 4629 2972
rect 4617 2941 4629 2944
rect 4663 2972 4675 2975
rect 4798 2972 4804 2984
rect 4663 2944 4804 2972
rect 4663 2941 4675 2944
rect 4617 2935 4675 2941
rect 4798 2932 4804 2944
rect 4856 2932 4862 2984
rect 4982 2932 4988 2984
rect 5040 2932 5046 2984
rect 5102 2975 5160 2981
rect 5102 2941 5114 2975
rect 5148 2972 5160 2975
rect 5626 2972 5632 2984
rect 5148 2944 5632 2972
rect 5148 2941 5160 2944
rect 5102 2935 5160 2941
rect 5626 2932 5632 2944
rect 5684 2932 5690 2984
rect 3605 2907 3663 2913
rect 3605 2873 3617 2907
rect 3651 2904 3663 2907
rect 4062 2904 4068 2916
rect 3651 2876 4068 2904
rect 3651 2873 3663 2876
rect 3605 2867 3663 2873
rect 4062 2864 4068 2876
rect 4120 2864 4126 2916
rect 1486 2796 1492 2848
rect 1544 2836 1550 2848
rect 2866 2836 2872 2848
rect 1544 2808 2872 2836
rect 1544 2796 1550 2808
rect 2866 2796 2872 2808
rect 2924 2796 2930 2848
rect 3970 2796 3976 2848
rect 4028 2836 4034 2848
rect 5736 2836 5764 3148
rect 7653 3145 7665 3148
rect 7699 3145 7711 3179
rect 7653 3139 7711 3145
rect 8110 3136 8116 3188
rect 8168 3176 8174 3188
rect 8389 3179 8447 3185
rect 8389 3176 8401 3179
rect 8168 3148 8401 3176
rect 8168 3136 8174 3148
rect 8389 3145 8401 3148
rect 8435 3145 8447 3179
rect 8389 3139 8447 3145
rect 9490 3136 9496 3188
rect 9548 3176 9554 3188
rect 11977 3179 12035 3185
rect 11977 3176 11989 3179
rect 9548 3148 11989 3176
rect 9548 3136 9554 3148
rect 11977 3145 11989 3148
rect 12023 3145 12035 3179
rect 11977 3139 12035 3145
rect 14182 3136 14188 3188
rect 14240 3176 14246 3188
rect 15013 3179 15071 3185
rect 15013 3176 15025 3179
rect 14240 3148 15025 3176
rect 14240 3136 14246 3148
rect 15013 3145 15025 3148
rect 15059 3145 15071 3179
rect 15013 3139 15071 3145
rect 15105 3179 15163 3185
rect 15105 3145 15117 3179
rect 15151 3176 15163 3179
rect 16206 3176 16212 3188
rect 15151 3148 16212 3176
rect 15151 3145 15163 3148
rect 15105 3139 15163 3145
rect 16206 3136 16212 3148
rect 16264 3176 16270 3188
rect 17221 3179 17279 3185
rect 16264 3148 16574 3176
rect 16264 3136 16270 3148
rect 6730 3108 6736 3120
rect 6656 3080 6736 3108
rect 5812 3043 5870 3049
rect 5812 3009 5824 3043
rect 5858 3009 5870 3043
rect 5812 3003 5870 3009
rect 5828 2972 5856 3003
rect 5902 3000 5908 3052
rect 5960 3000 5966 3052
rect 6656 3049 6684 3080
rect 6730 3068 6736 3080
rect 6788 3108 6794 3120
rect 6788 3080 8156 3108
rect 6788 3068 6794 3080
rect 6641 3043 6699 3049
rect 6641 3009 6653 3043
rect 6687 3009 6699 3043
rect 6641 3003 6699 3009
rect 7469 3043 7527 3049
rect 7469 3009 7481 3043
rect 7515 3040 7527 3043
rect 7558 3040 7564 3052
rect 7515 3012 7564 3040
rect 7515 3009 7527 3012
rect 7469 3003 7527 3009
rect 7558 3000 7564 3012
rect 7616 3000 7622 3052
rect 8128 3049 8156 3080
rect 9306 3068 9312 3120
rect 9364 3068 9370 3120
rect 11146 3108 11152 3120
rect 10534 3080 11152 3108
rect 11146 3068 11152 3080
rect 11204 3068 11210 3120
rect 14642 3108 14648 3120
rect 13740 3080 14648 3108
rect 7745 3043 7803 3049
rect 7745 3009 7757 3043
rect 7791 3009 7803 3043
rect 7745 3003 7803 3009
rect 8021 3043 8079 3049
rect 8021 3009 8033 3043
rect 8067 3009 8079 3043
rect 8021 3003 8079 3009
rect 8114 3043 8172 3049
rect 8114 3009 8126 3043
rect 8160 3009 8172 3043
rect 8114 3003 8172 3009
rect 5994 2972 6000 2984
rect 5828 2944 6000 2972
rect 5994 2932 6000 2944
rect 6052 2932 6058 2984
rect 6733 2975 6791 2981
rect 6733 2941 6745 2975
rect 6779 2972 6791 2975
rect 6779 2944 7328 2972
rect 6779 2941 6791 2944
rect 6733 2935 6791 2941
rect 7009 2907 7067 2913
rect 7009 2873 7021 2907
rect 7055 2904 7067 2907
rect 7190 2904 7196 2916
rect 7055 2876 7196 2904
rect 7055 2873 7067 2876
rect 7009 2867 7067 2873
rect 7190 2864 7196 2876
rect 7248 2864 7254 2916
rect 7300 2904 7328 2944
rect 7374 2932 7380 2984
rect 7432 2972 7438 2984
rect 7760 2972 7788 3003
rect 7432 2944 7788 2972
rect 8036 2972 8064 3003
rect 9030 3000 9036 3052
rect 9088 3000 9094 3052
rect 12069 3043 12127 3049
rect 12069 3009 12081 3043
rect 12115 3040 12127 3043
rect 12115 3012 12572 3040
rect 12115 3009 12127 3012
rect 12069 3003 12127 3009
rect 9398 2972 9404 2984
rect 8036 2944 9404 2972
rect 7432 2932 7438 2944
rect 8036 2904 8064 2944
rect 9398 2932 9404 2944
rect 9456 2932 9462 2984
rect 12161 2975 12219 2981
rect 12161 2941 12173 2975
rect 12207 2941 12219 2975
rect 12544 2972 12572 3012
rect 12618 3000 12624 3052
rect 12676 3000 12682 3052
rect 12805 3043 12863 3049
rect 12805 3009 12817 3043
rect 12851 3040 12863 3043
rect 12894 3040 12900 3052
rect 12851 3012 12900 3040
rect 12851 3009 12863 3012
rect 12805 3003 12863 3009
rect 12894 3000 12900 3012
rect 12952 3040 12958 3052
rect 13078 3040 13084 3052
rect 12952 3012 13084 3040
rect 12952 3000 12958 3012
rect 13078 3000 13084 3012
rect 13136 3000 13142 3052
rect 13740 3049 13768 3080
rect 14642 3068 14648 3080
rect 14700 3068 14706 3120
rect 16546 3108 16574 3148
rect 17221 3145 17233 3179
rect 17267 3176 17279 3179
rect 17586 3176 17592 3188
rect 17267 3148 17592 3176
rect 17267 3145 17279 3148
rect 17221 3139 17279 3145
rect 17586 3136 17592 3148
rect 17644 3136 17650 3188
rect 21542 3136 21548 3188
rect 21600 3136 21606 3188
rect 22002 3136 22008 3188
rect 22060 3136 22066 3188
rect 17313 3111 17371 3117
rect 17313 3108 17325 3111
rect 14936 3080 15792 3108
rect 16546 3080 17325 3108
rect 13725 3043 13783 3049
rect 13725 3009 13737 3043
rect 13771 3009 13783 3043
rect 13725 3003 13783 3009
rect 13814 3000 13820 3052
rect 13872 3040 13878 3052
rect 14185 3043 14243 3049
rect 14185 3040 14197 3043
rect 13872 3012 14197 3040
rect 13872 3000 13878 3012
rect 14185 3009 14197 3012
rect 14231 3009 14243 3043
rect 14185 3003 14243 3009
rect 14274 3000 14280 3052
rect 14332 3040 14338 3052
rect 14369 3043 14427 3049
rect 14369 3040 14381 3043
rect 14332 3012 14381 3040
rect 14332 3000 14338 3012
rect 14369 3009 14381 3012
rect 14415 3009 14427 3043
rect 14369 3003 14427 3009
rect 14936 2972 14964 3080
rect 15654 3040 15660 3052
rect 12544 2944 14964 2972
rect 15028 3012 15660 3040
rect 12161 2935 12219 2941
rect 7300 2876 8064 2904
rect 12066 2864 12072 2916
rect 12124 2904 12130 2916
rect 12176 2904 12204 2935
rect 12124 2876 12204 2904
rect 13909 2907 13967 2913
rect 12124 2864 12130 2876
rect 13909 2873 13921 2907
rect 13955 2904 13967 2907
rect 15028 2904 15056 3012
rect 15654 3000 15660 3012
rect 15712 3000 15718 3052
rect 15197 2975 15255 2981
rect 15197 2972 15209 2975
rect 13955 2876 15056 2904
rect 15120 2944 15209 2972
rect 13955 2873 13967 2876
rect 13909 2867 13967 2873
rect 4028 2808 5764 2836
rect 4028 2796 4034 2808
rect 7282 2796 7288 2848
rect 7340 2796 7346 2848
rect 9306 2796 9312 2848
rect 9364 2836 9370 2848
rect 10781 2839 10839 2845
rect 10781 2836 10793 2839
rect 9364 2808 10793 2836
rect 9364 2796 9370 2808
rect 10781 2805 10793 2808
rect 10827 2805 10839 2839
rect 10781 2799 10839 2805
rect 11238 2796 11244 2848
rect 11296 2836 11302 2848
rect 11609 2839 11667 2845
rect 11609 2836 11621 2839
rect 11296 2808 11621 2836
rect 11296 2796 11302 2808
rect 11609 2805 11621 2808
rect 11655 2805 11667 2839
rect 11609 2799 11667 2805
rect 12802 2796 12808 2848
rect 12860 2796 12866 2848
rect 14366 2796 14372 2848
rect 14424 2796 14430 2848
rect 14642 2796 14648 2848
rect 14700 2796 14706 2848
rect 14918 2796 14924 2848
rect 14976 2836 14982 2848
rect 15120 2836 15148 2944
rect 15197 2941 15209 2944
rect 15243 2941 15255 2975
rect 15197 2935 15255 2941
rect 15764 2904 15792 3080
rect 17313 3077 17325 3080
rect 17359 3077 17371 3111
rect 17313 3071 17371 3077
rect 21082 3068 21088 3120
rect 21140 3068 21146 3120
rect 15838 3000 15844 3052
rect 15896 3040 15902 3052
rect 16209 3043 16267 3049
rect 16209 3040 16221 3043
rect 15896 3012 16221 3040
rect 15896 3000 15902 3012
rect 16209 3009 16221 3012
rect 16255 3009 16267 3043
rect 16209 3003 16267 3009
rect 16393 3043 16451 3049
rect 16393 3009 16405 3043
rect 16439 3040 16451 3043
rect 16666 3040 16672 3052
rect 16439 3012 16672 3040
rect 16439 3009 16451 3012
rect 16393 3003 16451 3009
rect 16224 2972 16252 3003
rect 16666 3000 16672 3012
rect 16724 3040 16730 3052
rect 19702 3040 19708 3052
rect 16724 3012 19708 3040
rect 16724 3000 16730 3012
rect 19702 3000 19708 3012
rect 19760 3000 19766 3052
rect 19794 3000 19800 3052
rect 19852 3000 19858 3052
rect 21450 3000 21456 3052
rect 21508 3040 21514 3052
rect 21913 3043 21971 3049
rect 21913 3040 21925 3043
rect 21508 3012 21925 3040
rect 21508 3000 21514 3012
rect 21913 3009 21925 3012
rect 21959 3009 21971 3043
rect 21913 3003 21971 3009
rect 22097 3043 22155 3049
rect 22097 3009 22109 3043
rect 22143 3040 22155 3043
rect 23750 3040 23756 3052
rect 22143 3012 23756 3040
rect 22143 3009 22155 3012
rect 22097 3003 22155 3009
rect 23750 3000 23756 3012
rect 23808 3000 23814 3052
rect 16942 2972 16948 2984
rect 16224 2944 16948 2972
rect 16942 2932 16948 2944
rect 17000 2932 17006 2984
rect 17129 2975 17187 2981
rect 17129 2941 17141 2975
rect 17175 2941 17187 2975
rect 17129 2935 17187 2941
rect 15764 2876 16988 2904
rect 14976 2808 15148 2836
rect 16209 2839 16267 2845
rect 14976 2796 14982 2808
rect 16209 2805 16221 2839
rect 16255 2836 16267 2839
rect 16574 2836 16580 2848
rect 16255 2808 16580 2836
rect 16255 2805 16267 2808
rect 16209 2799 16267 2805
rect 16574 2796 16580 2808
rect 16632 2796 16638 2848
rect 16960 2836 16988 2876
rect 17034 2864 17040 2916
rect 17092 2904 17098 2916
rect 17144 2904 17172 2935
rect 17218 2932 17224 2984
rect 17276 2972 17282 2984
rect 19610 2972 19616 2984
rect 17276 2944 19616 2972
rect 17276 2932 17282 2944
rect 19610 2932 19616 2944
rect 19668 2932 19674 2984
rect 20070 2932 20076 2984
rect 20128 2932 20134 2984
rect 18506 2904 18512 2916
rect 17092 2876 17172 2904
rect 17604 2876 18512 2904
rect 17092 2864 17098 2876
rect 17604 2836 17632 2876
rect 18506 2864 18512 2876
rect 18564 2864 18570 2916
rect 16960 2808 17632 2836
rect 17681 2839 17739 2845
rect 17681 2805 17693 2839
rect 17727 2836 17739 2839
rect 18414 2836 18420 2848
rect 17727 2808 18420 2836
rect 17727 2805 17739 2808
rect 17681 2799 17739 2805
rect 18414 2796 18420 2808
rect 18472 2796 18478 2848
rect 1104 2746 25852 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 12214 2746
rect 12266 2694 12278 2746
rect 12330 2694 12342 2746
rect 12394 2694 12406 2746
rect 12458 2694 12470 2746
rect 12522 2694 20214 2746
rect 20266 2694 20278 2746
rect 20330 2694 20342 2746
rect 20394 2694 20406 2746
rect 20458 2694 20470 2746
rect 20522 2694 25852 2746
rect 1104 2672 25852 2694
rect 8481 2635 8539 2641
rect 8481 2601 8493 2635
rect 8527 2632 8539 2635
rect 8570 2632 8576 2644
rect 8527 2604 8576 2632
rect 8527 2601 8539 2604
rect 8481 2595 8539 2601
rect 8570 2592 8576 2604
rect 8628 2592 8634 2644
rect 12618 2592 12624 2644
rect 12676 2632 12682 2644
rect 13722 2632 13728 2644
rect 12676 2604 13728 2632
rect 12676 2592 12682 2604
rect 2866 2456 2872 2508
rect 2924 2496 2930 2508
rect 3881 2499 3939 2505
rect 3881 2496 3893 2499
rect 2924 2468 3893 2496
rect 2924 2456 2930 2468
rect 3881 2465 3893 2468
rect 3927 2465 3939 2499
rect 3881 2459 3939 2465
rect 5629 2499 5687 2505
rect 5629 2465 5641 2499
rect 5675 2465 5687 2499
rect 5629 2459 5687 2465
rect 3513 2431 3571 2437
rect 3513 2397 3525 2431
rect 3559 2397 3571 2431
rect 5644 2428 5672 2459
rect 7006 2456 7012 2508
rect 7064 2456 7070 2508
rect 7190 2456 7196 2508
rect 7248 2496 7254 2508
rect 7653 2499 7711 2505
rect 7653 2496 7665 2499
rect 7248 2468 7665 2496
rect 7248 2456 7254 2468
rect 7653 2465 7665 2468
rect 7699 2496 7711 2499
rect 7699 2468 8432 2496
rect 7699 2465 7711 2468
rect 7653 2459 7711 2465
rect 5905 2431 5963 2437
rect 5905 2428 5917 2431
rect 5644 2400 5917 2428
rect 3513 2391 3571 2397
rect 5905 2397 5917 2400
rect 5951 2428 5963 2431
rect 5994 2428 6000 2440
rect 5951 2400 6000 2428
rect 5951 2397 5963 2400
rect 5905 2391 5963 2397
rect 3142 2252 3148 2304
rect 3200 2292 3206 2304
rect 3329 2295 3387 2301
rect 3329 2292 3341 2295
rect 3200 2264 3341 2292
rect 3200 2252 3206 2264
rect 3329 2261 3341 2264
rect 3375 2261 3387 2295
rect 3528 2292 3556 2391
rect 5994 2388 6000 2400
rect 6052 2388 6058 2440
rect 6089 2431 6147 2437
rect 6089 2397 6101 2431
rect 6135 2428 6147 2431
rect 7466 2428 7472 2440
rect 6135 2400 7472 2428
rect 6135 2397 6147 2400
rect 6089 2391 6147 2397
rect 7466 2388 7472 2400
rect 7524 2388 7530 2440
rect 8404 2437 8432 2468
rect 9858 2456 9864 2508
rect 9916 2496 9922 2508
rect 10870 2496 10876 2508
rect 9916 2468 10876 2496
rect 9916 2456 9922 2468
rect 10870 2456 10876 2468
rect 10928 2456 10934 2508
rect 7745 2431 7803 2437
rect 7745 2397 7757 2431
rect 7791 2397 7803 2431
rect 7745 2391 7803 2397
rect 8389 2431 8447 2437
rect 8389 2397 8401 2431
rect 8435 2397 8447 2431
rect 8389 2391 8447 2397
rect 8573 2431 8631 2437
rect 8573 2397 8585 2431
rect 8619 2428 8631 2431
rect 9122 2428 9128 2440
rect 8619 2400 9128 2428
rect 8619 2397 8631 2400
rect 8573 2391 8631 2397
rect 4157 2363 4215 2369
rect 4157 2329 4169 2363
rect 4203 2360 4215 2363
rect 4430 2360 4436 2372
rect 4203 2332 4436 2360
rect 4203 2329 4215 2332
rect 4157 2323 4215 2329
rect 4430 2320 4436 2332
rect 4488 2320 4494 2372
rect 4614 2320 4620 2372
rect 4672 2320 4678 2372
rect 5460 2332 6408 2360
rect 5460 2292 5488 2332
rect 3528 2264 5488 2292
rect 5997 2295 6055 2301
rect 3329 2255 3387 2261
rect 5997 2261 6009 2295
rect 6043 2292 6055 2295
rect 6270 2292 6276 2304
rect 6043 2264 6276 2292
rect 6043 2261 6055 2264
rect 5997 2255 6055 2261
rect 6270 2252 6276 2264
rect 6328 2252 6334 2304
rect 6380 2301 6408 2332
rect 6454 2320 6460 2372
rect 6512 2360 6518 2372
rect 6730 2360 6736 2372
rect 6512 2332 6736 2360
rect 6512 2320 6518 2332
rect 6730 2320 6736 2332
rect 6788 2320 6794 2372
rect 7760 2360 7788 2391
rect 8588 2360 8616 2391
rect 9122 2388 9128 2400
rect 9180 2388 9186 2440
rect 13078 2388 13084 2440
rect 13136 2428 13142 2440
rect 13188 2437 13216 2604
rect 13722 2592 13728 2604
rect 13780 2592 13786 2644
rect 14182 2592 14188 2644
rect 14240 2592 14246 2644
rect 16206 2592 16212 2644
rect 16264 2592 16270 2644
rect 13906 2496 13912 2508
rect 13372 2468 13912 2496
rect 13372 2437 13400 2468
rect 13173 2431 13231 2437
rect 13173 2428 13185 2431
rect 13136 2400 13185 2428
rect 13136 2388 13142 2400
rect 13173 2397 13185 2400
rect 13219 2397 13231 2431
rect 13173 2391 13231 2397
rect 13357 2431 13415 2437
rect 13357 2397 13369 2431
rect 13403 2397 13415 2431
rect 13357 2391 13415 2397
rect 13633 2431 13691 2437
rect 13633 2397 13645 2431
rect 13679 2428 13691 2431
rect 13722 2428 13728 2440
rect 13679 2400 13728 2428
rect 13679 2397 13691 2400
rect 13633 2391 13691 2397
rect 13722 2388 13728 2400
rect 13780 2388 13786 2440
rect 13832 2437 13860 2468
rect 13906 2456 13912 2468
rect 13964 2496 13970 2508
rect 14274 2496 14280 2508
rect 13964 2468 14280 2496
rect 13964 2456 13970 2468
rect 14274 2456 14280 2468
rect 14332 2456 14338 2508
rect 15654 2456 15660 2508
rect 15712 2456 15718 2508
rect 15930 2456 15936 2508
rect 15988 2496 15994 2508
rect 16666 2496 16672 2508
rect 15988 2468 16672 2496
rect 15988 2456 15994 2468
rect 16666 2456 16672 2468
rect 16724 2456 16730 2508
rect 19797 2499 19855 2505
rect 19797 2465 19809 2499
rect 19843 2496 19855 2499
rect 19886 2496 19892 2508
rect 19843 2468 19892 2496
rect 19843 2465 19855 2468
rect 19797 2459 19855 2465
rect 19886 2456 19892 2468
rect 19944 2456 19950 2508
rect 19978 2456 19984 2508
rect 20036 2456 20042 2508
rect 13817 2431 13875 2437
rect 13817 2397 13829 2431
rect 13863 2397 13875 2431
rect 13817 2391 13875 2397
rect 16574 2388 16580 2440
rect 16632 2388 16638 2440
rect 17957 2431 18015 2437
rect 17957 2397 17969 2431
rect 18003 2397 18015 2431
rect 17957 2391 18015 2397
rect 7760 2332 8616 2360
rect 11146 2320 11152 2372
rect 11204 2320 11210 2372
rect 12802 2360 12808 2372
rect 12374 2332 12808 2360
rect 12802 2320 12808 2332
rect 12860 2320 12866 2372
rect 13265 2363 13323 2369
rect 13265 2329 13277 2363
rect 13311 2360 13323 2363
rect 17681 2363 17739 2369
rect 13311 2332 14490 2360
rect 13311 2329 13323 2332
rect 13265 2323 13323 2329
rect 17681 2329 17693 2363
rect 17727 2329 17739 2363
rect 17681 2323 17739 2329
rect 6365 2295 6423 2301
rect 6365 2261 6377 2295
rect 6411 2261 6423 2295
rect 6365 2255 6423 2261
rect 6822 2252 6828 2304
rect 6880 2252 6886 2304
rect 8110 2252 8116 2304
rect 8168 2252 8174 2304
rect 12158 2252 12164 2304
rect 12216 2292 12222 2304
rect 12621 2295 12679 2301
rect 12621 2292 12633 2295
rect 12216 2264 12633 2292
rect 12216 2252 12222 2264
rect 12621 2261 12633 2264
rect 12667 2261 12679 2295
rect 12621 2255 12679 2261
rect 13725 2295 13783 2301
rect 13725 2261 13737 2295
rect 13771 2292 13783 2295
rect 17494 2292 17500 2304
rect 13771 2264 17500 2292
rect 13771 2261 13783 2264
rect 13725 2255 13783 2261
rect 17494 2252 17500 2264
rect 17552 2252 17558 2304
rect 17696 2292 17724 2323
rect 17770 2320 17776 2372
rect 17828 2360 17834 2372
rect 17972 2360 18000 2391
rect 18414 2388 18420 2440
rect 18472 2388 18478 2440
rect 18785 2431 18843 2437
rect 18785 2397 18797 2431
rect 18831 2428 18843 2431
rect 18831 2400 19380 2428
rect 18831 2397 18843 2400
rect 18785 2391 18843 2397
rect 17828 2332 18000 2360
rect 17828 2320 17834 2332
rect 18233 2295 18291 2301
rect 18233 2292 18245 2295
rect 17696 2264 18245 2292
rect 18233 2261 18245 2264
rect 18279 2261 18291 2295
rect 18233 2255 18291 2261
rect 18969 2295 19027 2301
rect 18969 2261 18981 2295
rect 19015 2292 19027 2295
rect 19058 2292 19064 2304
rect 19015 2264 19064 2292
rect 19015 2261 19027 2264
rect 18969 2255 19027 2261
rect 19058 2252 19064 2264
rect 19116 2252 19122 2304
rect 19352 2301 19380 2400
rect 19610 2388 19616 2440
rect 19668 2428 19674 2440
rect 20349 2431 20407 2437
rect 20349 2428 20361 2431
rect 19668 2400 20361 2428
rect 19668 2388 19674 2400
rect 20349 2397 20361 2400
rect 20395 2397 20407 2431
rect 20349 2391 20407 2397
rect 20533 2431 20591 2437
rect 20533 2397 20545 2431
rect 20579 2428 20591 2431
rect 20622 2428 20628 2440
rect 20579 2400 20628 2428
rect 20579 2397 20591 2400
rect 20533 2391 20591 2397
rect 20622 2388 20628 2400
rect 20680 2388 20686 2440
rect 19337 2295 19395 2301
rect 19337 2261 19349 2295
rect 19383 2261 19395 2295
rect 19337 2255 19395 2261
rect 19702 2252 19708 2304
rect 19760 2252 19766 2304
rect 20438 2252 20444 2304
rect 20496 2252 20502 2304
rect 1104 2202 25852 2224
rect 1104 2150 8214 2202
rect 8266 2150 8278 2202
rect 8330 2150 8342 2202
rect 8394 2150 8406 2202
rect 8458 2150 8470 2202
rect 8522 2150 16214 2202
rect 16266 2150 16278 2202
rect 16330 2150 16342 2202
rect 16394 2150 16406 2202
rect 16458 2150 16470 2202
rect 16522 2150 24214 2202
rect 24266 2150 24278 2202
rect 24330 2150 24342 2202
rect 24394 2150 24406 2202
rect 24458 2150 24470 2202
rect 24522 2150 25852 2202
rect 1104 2128 25852 2150
rect 4890 2048 4896 2100
rect 4948 2048 4954 2100
rect 5626 2048 5632 2100
rect 5684 2048 5690 2100
rect 7193 2091 7251 2097
rect 7193 2057 7205 2091
rect 7239 2088 7251 2091
rect 7742 2088 7748 2100
rect 7239 2060 7748 2088
rect 7239 2057 7251 2060
rect 7193 2051 7251 2057
rect 7742 2048 7748 2060
rect 7800 2048 7806 2100
rect 9490 2048 9496 2100
rect 9548 2048 9554 2100
rect 10796 2060 11376 2088
rect 3142 1980 3148 2032
rect 3200 1980 3206 2032
rect 4154 1980 4160 2032
rect 4212 1980 4218 2032
rect 4430 1980 4436 2032
rect 4488 2020 4494 2032
rect 6457 2023 6515 2029
rect 6457 2020 6469 2023
rect 4488 1992 6469 2020
rect 4488 1980 4494 1992
rect 6457 1989 6469 1992
rect 6503 1989 6515 2023
rect 10796 2020 10824 2060
rect 6457 1983 6515 1989
rect 6564 1992 7604 2020
rect 10534 1992 10824 2020
rect 2866 1912 2872 1964
rect 2924 1912 2930 1964
rect 5902 1952 5908 1964
rect 5863 1924 5908 1952
rect 5902 1912 5908 1924
rect 5960 1912 5966 1964
rect 5994 1912 6000 1964
rect 6052 1952 6058 1964
rect 6564 1952 6592 1992
rect 7576 1964 7604 1992
rect 10870 1980 10876 2032
rect 10928 2020 10934 2032
rect 11348 2020 11376 2060
rect 12158 2048 12164 2100
rect 12216 2088 12222 2100
rect 12253 2091 12311 2097
rect 12253 2088 12265 2091
rect 12216 2060 12265 2088
rect 12216 2048 12222 2060
rect 12253 2057 12265 2060
rect 12299 2057 12311 2091
rect 12253 2051 12311 2057
rect 12345 2091 12403 2097
rect 12345 2057 12357 2091
rect 12391 2088 12403 2091
rect 13541 2091 13599 2097
rect 13541 2088 13553 2091
rect 12391 2060 13553 2088
rect 12391 2057 12403 2060
rect 12345 2051 12403 2057
rect 13541 2057 13553 2060
rect 13587 2057 13599 2091
rect 13541 2051 13599 2057
rect 16666 2048 16672 2100
rect 16724 2088 16730 2100
rect 17770 2088 17776 2100
rect 16724 2060 17776 2088
rect 16724 2048 16730 2060
rect 12989 2023 13047 2029
rect 12989 2020 13001 2023
rect 10928 1992 11284 2020
rect 11348 1992 13001 2020
rect 10928 1980 10934 1992
rect 6052 1924 6592 1952
rect 6641 1955 6699 1961
rect 6052 1912 6058 1924
rect 6641 1921 6653 1955
rect 6687 1952 6699 1955
rect 7282 1952 7288 1964
rect 6687 1924 7288 1952
rect 6687 1921 6699 1924
rect 6641 1915 6699 1921
rect 7282 1912 7288 1924
rect 7340 1912 7346 1964
rect 7558 1912 7564 1964
rect 7616 1912 7622 1964
rect 8662 1912 8668 1964
rect 8720 1912 8726 1964
rect 11256 1961 11284 1992
rect 12989 1989 13001 1992
rect 13035 1989 13047 2023
rect 12989 1983 13047 1989
rect 14366 1980 14372 2032
rect 14424 1980 14430 2032
rect 15010 1980 15016 2032
rect 15068 1980 15074 2032
rect 11241 1955 11299 1961
rect 11241 1921 11253 1955
rect 11287 1921 11299 1955
rect 11241 1915 11299 1921
rect 12066 1912 12072 1964
rect 12124 1912 12130 1964
rect 12894 1912 12900 1964
rect 12952 1912 12958 1964
rect 13078 1912 13084 1964
rect 13136 1912 13142 1964
rect 16776 1961 16804 2060
rect 17770 2048 17776 2060
rect 17828 2048 17834 2100
rect 18506 2048 18512 2100
rect 18564 2048 18570 2100
rect 17494 1980 17500 2032
rect 17552 1980 17558 2032
rect 19058 1980 19064 2032
rect 19116 1980 19122 2032
rect 20438 2020 20444 2032
rect 20286 1992 20444 2020
rect 20438 1980 20444 1992
rect 20496 1980 20502 2032
rect 15289 1955 15347 1961
rect 15289 1921 15301 1955
rect 15335 1952 15347 1955
rect 16761 1955 16819 1961
rect 16761 1952 16773 1955
rect 15335 1924 16773 1952
rect 15335 1921 15347 1924
rect 15289 1915 15347 1921
rect 16761 1921 16773 1924
rect 16807 1921 16819 1955
rect 16761 1915 16819 1921
rect 4617 1887 4675 1893
rect 4617 1853 4629 1887
rect 4663 1884 4675 1887
rect 4890 1884 4896 1896
rect 4663 1856 4896 1884
rect 4663 1853 4675 1856
rect 4617 1847 4675 1853
rect 4890 1844 4896 1856
rect 4948 1884 4954 1896
rect 5353 1887 5411 1893
rect 5353 1884 5365 1887
rect 4948 1856 5365 1884
rect 4948 1844 4954 1856
rect 5353 1853 5365 1856
rect 5399 1853 5411 1887
rect 5353 1847 5411 1853
rect 5074 1776 5080 1828
rect 5132 1776 5138 1828
rect 5368 1816 5396 1847
rect 6270 1844 6276 1896
rect 6328 1884 6334 1896
rect 6730 1884 6736 1896
rect 6328 1856 6736 1884
rect 6328 1844 6334 1856
rect 6730 1844 6736 1856
rect 6788 1884 6794 1896
rect 6825 1887 6883 1893
rect 6825 1884 6837 1887
rect 6788 1856 6837 1884
rect 6788 1844 6794 1856
rect 6825 1853 6837 1856
rect 6871 1853 6883 1887
rect 6825 1847 6883 1853
rect 6917 1887 6975 1893
rect 6917 1853 6929 1887
rect 6963 1853 6975 1887
rect 6917 1847 6975 1853
rect 6454 1816 6460 1828
rect 5368 1788 6460 1816
rect 6454 1776 6460 1788
rect 6512 1776 6518 1828
rect 6932 1748 6960 1847
rect 7374 1844 7380 1896
rect 7432 1844 7438 1896
rect 7466 1844 7472 1896
rect 7524 1844 7530 1896
rect 7653 1887 7711 1893
rect 7653 1853 7665 1887
rect 7699 1884 7711 1887
rect 8386 1884 8392 1896
rect 7699 1856 8392 1884
rect 7699 1853 7711 1856
rect 7653 1847 7711 1853
rect 8386 1844 8392 1856
rect 8444 1844 8450 1896
rect 8757 1887 8815 1893
rect 8757 1853 8769 1887
rect 8803 1884 8815 1887
rect 9214 1884 9220 1896
rect 8803 1856 9220 1884
rect 8803 1853 8815 1856
rect 8757 1847 8815 1853
rect 9214 1844 9220 1856
rect 9272 1844 9278 1896
rect 10962 1844 10968 1896
rect 11020 1844 11026 1896
rect 12084 1884 12112 1912
rect 12437 1887 12495 1893
rect 12437 1884 12449 1887
rect 12084 1856 12449 1884
rect 12437 1853 12449 1856
rect 12483 1853 12495 1887
rect 12437 1847 12495 1853
rect 17034 1844 17040 1896
rect 17092 1844 17098 1896
rect 17770 1844 17776 1896
rect 17828 1884 17834 1896
rect 18785 1887 18843 1893
rect 18785 1884 18797 1887
rect 17828 1856 18797 1884
rect 17828 1844 17834 1856
rect 18785 1853 18797 1856
rect 18831 1853 18843 1887
rect 18785 1847 18843 1853
rect 7484 1816 7512 1844
rect 8297 1819 8355 1825
rect 8297 1816 8309 1819
rect 7484 1788 8309 1816
rect 8297 1785 8309 1788
rect 8343 1785 8355 1819
rect 8297 1779 8355 1785
rect 8846 1748 8852 1760
rect 6932 1720 8852 1748
rect 8846 1708 8852 1720
rect 8904 1708 8910 1760
rect 11790 1708 11796 1760
rect 11848 1748 11854 1760
rect 11885 1751 11943 1757
rect 11885 1748 11897 1751
rect 11848 1720 11897 1748
rect 11848 1708 11854 1720
rect 11885 1717 11897 1720
rect 11931 1717 11943 1751
rect 11885 1711 11943 1717
rect 13538 1708 13544 1760
rect 13596 1708 13602 1760
rect 19702 1708 19708 1760
rect 19760 1748 19766 1760
rect 20533 1751 20591 1757
rect 20533 1748 20545 1751
rect 19760 1720 20545 1748
rect 19760 1708 19766 1720
rect 20533 1717 20545 1720
rect 20579 1717 20591 1751
rect 20533 1711 20591 1717
rect 1104 1658 25852 1680
rect 1104 1606 4214 1658
rect 4266 1606 4278 1658
rect 4330 1606 4342 1658
rect 4394 1606 4406 1658
rect 4458 1606 4470 1658
rect 4522 1606 12214 1658
rect 12266 1606 12278 1658
rect 12330 1606 12342 1658
rect 12394 1606 12406 1658
rect 12458 1606 12470 1658
rect 12522 1606 20214 1658
rect 20266 1606 20278 1658
rect 20330 1606 20342 1658
rect 20394 1606 20406 1658
rect 20458 1606 20470 1658
rect 20522 1606 25852 1658
rect 1104 1584 25852 1606
rect 4801 1547 4859 1553
rect 4801 1513 4813 1547
rect 4847 1544 4859 1547
rect 4982 1544 4988 1556
rect 4847 1516 4988 1544
rect 4847 1513 4859 1516
rect 4801 1507 4859 1513
rect 4982 1504 4988 1516
rect 5040 1504 5046 1556
rect 6822 1504 6828 1556
rect 6880 1504 6886 1556
rect 8386 1504 8392 1556
rect 8444 1504 8450 1556
rect 10962 1504 10968 1556
rect 11020 1544 11026 1556
rect 11057 1547 11115 1553
rect 11057 1544 11069 1547
rect 11020 1516 11069 1544
rect 11020 1504 11026 1516
rect 11057 1513 11069 1516
rect 11103 1513 11115 1547
rect 11057 1507 11115 1513
rect 11146 1504 11152 1556
rect 11204 1544 11210 1556
rect 11609 1547 11667 1553
rect 11609 1544 11621 1547
rect 11204 1516 11621 1544
rect 11204 1504 11210 1516
rect 11609 1513 11621 1516
rect 11655 1513 11667 1547
rect 11609 1507 11667 1513
rect 17034 1504 17040 1556
rect 17092 1504 17098 1556
rect 8662 1436 8668 1488
rect 8720 1476 8726 1488
rect 9217 1479 9275 1485
rect 9217 1476 9229 1479
rect 8720 1448 9229 1476
rect 8720 1436 8726 1448
rect 9217 1445 9229 1448
rect 9263 1476 9275 1479
rect 12066 1476 12072 1488
rect 9263 1448 12072 1476
rect 9263 1445 9275 1448
rect 9217 1439 9275 1445
rect 12066 1436 12072 1448
rect 12124 1436 12130 1488
rect 14918 1436 14924 1488
rect 14976 1436 14982 1488
rect 842 1368 848 1420
rect 900 1408 906 1420
rect 1489 1411 1547 1417
rect 1489 1408 1501 1411
rect 900 1380 1501 1408
rect 900 1368 906 1380
rect 1489 1377 1501 1380
rect 1535 1377 1547 1411
rect 1489 1371 1547 1377
rect 7193 1411 7251 1417
rect 7193 1377 7205 1411
rect 7239 1408 7251 1411
rect 7374 1408 7380 1420
rect 7239 1380 7380 1408
rect 7239 1377 7251 1380
rect 7193 1371 7251 1377
rect 7374 1368 7380 1380
rect 7432 1408 7438 1420
rect 7561 1411 7619 1417
rect 7561 1408 7573 1411
rect 7432 1380 7573 1408
rect 7432 1368 7438 1380
rect 7561 1377 7573 1380
rect 7607 1377 7619 1411
rect 7561 1371 7619 1377
rect 8021 1411 8079 1417
rect 8021 1377 8033 1411
rect 8067 1408 8079 1411
rect 8110 1408 8116 1420
rect 8067 1380 8116 1408
rect 8067 1377 8079 1380
rect 8021 1371 8079 1377
rect 8110 1368 8116 1380
rect 8168 1368 8174 1420
rect 14936 1408 14964 1436
rect 15105 1411 15163 1417
rect 15105 1408 15117 1411
rect 14936 1380 15117 1408
rect 15105 1377 15117 1380
rect 15151 1408 15163 1411
rect 18141 1411 18199 1417
rect 18141 1408 18153 1411
rect 15151 1380 18153 1408
rect 15151 1377 15163 1380
rect 15105 1371 15163 1377
rect 18141 1377 18153 1380
rect 18187 1377 18199 1411
rect 19702 1408 19708 1420
rect 18141 1371 18199 1377
rect 18616 1380 19708 1408
rect 2866 1300 2872 1352
rect 2924 1340 2930 1352
rect 3237 1343 3295 1349
rect 3237 1340 3249 1343
rect 2924 1312 3249 1340
rect 2924 1300 2930 1312
rect 3237 1309 3249 1312
rect 3283 1309 3295 1343
rect 4890 1340 4896 1352
rect 4851 1312 4896 1340
rect 3237 1303 3295 1309
rect 4890 1300 4896 1312
rect 4948 1300 4954 1352
rect 4985 1343 5043 1349
rect 4985 1309 4997 1343
rect 5031 1340 5043 1343
rect 5074 1340 5080 1352
rect 5031 1312 5080 1340
rect 5031 1309 5043 1312
rect 4985 1303 5043 1309
rect 5074 1300 5080 1312
rect 5132 1300 5138 1352
rect 6730 1300 6736 1352
rect 6788 1340 6794 1352
rect 7101 1343 7159 1349
rect 7101 1340 7113 1343
rect 6788 1312 7113 1340
rect 6788 1300 6794 1312
rect 7101 1309 7113 1312
rect 7147 1309 7159 1343
rect 7101 1303 7159 1309
rect 7929 1343 7987 1349
rect 7929 1309 7941 1343
rect 7975 1309 7987 1343
rect 8128 1340 8156 1368
rect 8389 1343 8447 1349
rect 8389 1340 8401 1343
rect 8128 1312 8401 1340
rect 7929 1303 7987 1309
rect 8389 1309 8401 1312
rect 8435 1309 8447 1343
rect 8389 1303 8447 1309
rect 8573 1343 8631 1349
rect 8573 1309 8585 1343
rect 8619 1340 8631 1343
rect 8619 1312 9076 1340
rect 8619 1309 8631 1312
rect 8573 1303 8631 1309
rect 7944 1272 7972 1303
rect 8588 1272 8616 1303
rect 7944 1244 8616 1272
rect 9048 1213 9076 1312
rect 9214 1300 9220 1352
rect 9272 1340 9278 1352
rect 9493 1343 9551 1349
rect 9493 1340 9505 1343
rect 9272 1312 9505 1340
rect 9272 1300 9278 1312
rect 9493 1309 9505 1312
rect 9539 1309 9551 1343
rect 9493 1303 9551 1309
rect 11238 1300 11244 1352
rect 11296 1300 11302 1352
rect 11790 1300 11796 1352
rect 11848 1300 11854 1352
rect 13538 1300 13544 1352
rect 13596 1340 13602 1352
rect 14921 1343 14979 1349
rect 14921 1340 14933 1343
rect 13596 1312 14933 1340
rect 13596 1300 13602 1312
rect 14921 1309 14933 1312
rect 14967 1309 14979 1343
rect 14921 1303 14979 1309
rect 17221 1343 17279 1349
rect 17221 1309 17233 1343
rect 17267 1340 17279 1343
rect 17957 1343 18015 1349
rect 17267 1312 17632 1340
rect 17267 1309 17279 1312
rect 17221 1303 17279 1309
rect 15013 1275 15071 1281
rect 15013 1241 15025 1275
rect 15059 1272 15071 1275
rect 15102 1272 15108 1284
rect 15059 1244 15108 1272
rect 15059 1241 15071 1244
rect 15013 1235 15071 1241
rect 15102 1232 15108 1244
rect 15160 1232 15166 1284
rect 9033 1207 9091 1213
rect 9033 1173 9045 1207
rect 9079 1173 9091 1207
rect 9033 1167 9091 1173
rect 14550 1164 14556 1216
rect 14608 1164 14614 1216
rect 17604 1213 17632 1312
rect 17957 1309 17969 1343
rect 18003 1340 18015 1343
rect 18506 1340 18512 1352
rect 18003 1312 18512 1340
rect 18003 1309 18015 1312
rect 17957 1303 18015 1309
rect 18506 1300 18512 1312
rect 18564 1300 18570 1352
rect 18049 1275 18107 1281
rect 18049 1241 18061 1275
rect 18095 1272 18107 1275
rect 18616 1272 18644 1380
rect 19702 1368 19708 1380
rect 19760 1368 19766 1420
rect 18095 1244 18644 1272
rect 18095 1241 18107 1244
rect 18049 1235 18107 1241
rect 17589 1207 17647 1213
rect 17589 1173 17601 1207
rect 17635 1173 17647 1207
rect 17589 1167 17647 1173
rect 1104 1114 25852 1136
rect 1104 1062 8214 1114
rect 8266 1062 8278 1114
rect 8330 1062 8342 1114
rect 8394 1062 8406 1114
rect 8458 1062 8470 1114
rect 8522 1062 16214 1114
rect 16266 1062 16278 1114
rect 16330 1062 16342 1114
rect 16394 1062 16406 1114
rect 16458 1062 16470 1114
rect 16522 1062 24214 1114
rect 24266 1062 24278 1114
rect 24330 1062 24342 1114
rect 24394 1062 24406 1114
rect 24458 1062 24470 1114
rect 24522 1062 25852 1114
rect 1104 1040 25852 1062
<< via1 >>
rect 1400 21292 1452 21344
rect 13176 21292 13228 21344
rect 3608 21224 3660 21276
rect 14556 21224 14608 21276
rect 5356 21156 5408 21208
rect 14280 21156 14332 21208
rect 9128 20952 9180 21004
rect 9956 20952 10008 21004
rect 15568 20952 15620 21004
rect 7380 20884 7432 20936
rect 15292 20884 15344 20936
rect 9404 20816 9456 20868
rect 14648 20816 14700 20868
rect 11428 20748 11480 20800
rect 14096 20748 14148 20800
rect 8214 20646 8266 20698
rect 8278 20646 8330 20698
rect 8342 20646 8394 20698
rect 8406 20646 8458 20698
rect 8470 20646 8522 20698
rect 16214 20646 16266 20698
rect 16278 20646 16330 20698
rect 16342 20646 16394 20698
rect 16406 20646 16458 20698
rect 16470 20646 16522 20698
rect 24214 20646 24266 20698
rect 24278 20646 24330 20698
rect 24342 20646 24394 20698
rect 24406 20646 24458 20698
rect 24470 20646 24522 20698
rect 4712 20408 4764 20460
rect 4896 20408 4948 20460
rect 8760 20544 8812 20596
rect 9864 20476 9916 20528
rect 7380 20451 7432 20460
rect 7380 20417 7389 20451
rect 7389 20417 7423 20451
rect 7423 20417 7432 20451
rect 7380 20408 7432 20417
rect 8576 20408 8628 20460
rect 9128 20451 9180 20460
rect 9128 20417 9137 20451
rect 9137 20417 9171 20451
rect 9171 20417 9180 20451
rect 9128 20408 9180 20417
rect 9312 20408 9364 20460
rect 11980 20476 12032 20528
rect 13728 20408 13780 20460
rect 16304 20544 16356 20596
rect 15476 20408 15528 20460
rect 204 20340 256 20392
rect 5172 20383 5224 20392
rect 5172 20349 5181 20383
rect 5181 20349 5215 20383
rect 5215 20349 5224 20383
rect 5172 20340 5224 20349
rect 10048 20340 10100 20392
rect 11152 20340 11204 20392
rect 11244 20340 11296 20392
rect 12716 20340 12768 20392
rect 13636 20340 13688 20392
rect 15660 20340 15712 20392
rect 15752 20383 15804 20392
rect 15752 20349 15761 20383
rect 15761 20349 15795 20383
rect 15795 20349 15804 20383
rect 15752 20340 15804 20349
rect 10232 20272 10284 20324
rect 12072 20315 12124 20324
rect 12072 20281 12081 20315
rect 12081 20281 12115 20315
rect 12115 20281 12124 20315
rect 12072 20272 12124 20281
rect 14188 20315 14240 20324
rect 14188 20281 14197 20315
rect 14197 20281 14231 20315
rect 14231 20281 14240 20315
rect 14188 20272 14240 20281
rect 17224 20272 17276 20324
rect 5356 20247 5408 20256
rect 5356 20213 5365 20247
rect 5365 20213 5399 20247
rect 5399 20213 5408 20247
rect 5356 20204 5408 20213
rect 5540 20204 5592 20256
rect 5908 20204 5960 20256
rect 7472 20204 7524 20256
rect 9404 20204 9456 20256
rect 9496 20204 9548 20256
rect 12716 20247 12768 20256
rect 12716 20213 12725 20247
rect 12725 20213 12759 20247
rect 12759 20213 12768 20247
rect 12716 20204 12768 20213
rect 15016 20247 15068 20256
rect 15016 20213 15025 20247
rect 15025 20213 15059 20247
rect 15059 20213 15068 20247
rect 15016 20204 15068 20213
rect 15200 20204 15252 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 12214 20102 12266 20154
rect 12278 20102 12330 20154
rect 12342 20102 12394 20154
rect 12406 20102 12458 20154
rect 12470 20102 12522 20154
rect 20214 20102 20266 20154
rect 20278 20102 20330 20154
rect 20342 20102 20394 20154
rect 20406 20102 20458 20154
rect 20470 20102 20522 20154
rect 9404 19975 9456 19984
rect 9404 19941 9413 19975
rect 9413 19941 9447 19975
rect 9447 19941 9456 19975
rect 9404 19932 9456 19941
rect 9864 20043 9916 20052
rect 9864 20009 9873 20043
rect 9873 20009 9907 20043
rect 9907 20009 9916 20043
rect 9864 20000 9916 20009
rect 11980 20000 12032 20052
rect 12072 20000 12124 20052
rect 5908 19864 5960 19916
rect 4896 19796 4948 19848
rect 5448 19796 5500 19848
rect 7012 19796 7064 19848
rect 9496 19864 9548 19916
rect 10048 19907 10100 19916
rect 10048 19873 10057 19907
rect 10057 19873 10091 19907
rect 10091 19873 10100 19907
rect 10048 19864 10100 19873
rect 10232 19864 10284 19916
rect 11152 19975 11204 19984
rect 11152 19941 11161 19975
rect 11161 19941 11195 19975
rect 11195 19941 11204 19975
rect 11152 19932 11204 19941
rect 13452 20000 13504 20052
rect 14188 20043 14240 20052
rect 14188 20009 14197 20043
rect 14197 20009 14231 20043
rect 14231 20009 14240 20043
rect 14188 20000 14240 20009
rect 10416 19864 10468 19916
rect 13728 19975 13780 19984
rect 13728 19941 13737 19975
rect 13737 19941 13771 19975
rect 13771 19941 13780 19975
rect 13728 19932 13780 19941
rect 15384 20000 15436 20052
rect 15476 20043 15528 20052
rect 15476 20009 15485 20043
rect 15485 20009 15519 20043
rect 15519 20009 15528 20043
rect 15476 20000 15528 20009
rect 16304 20043 16356 20052
rect 16304 20009 16313 20043
rect 16313 20009 16347 20043
rect 16347 20009 16356 20043
rect 16304 20000 16356 20009
rect 17224 20043 17276 20052
rect 17224 20009 17233 20043
rect 17233 20009 17267 20043
rect 17267 20009 17276 20043
rect 17224 20000 17276 20009
rect 15016 19932 15068 19984
rect 8944 19796 8996 19848
rect 9128 19796 9180 19848
rect 7380 19728 7432 19780
rect 11612 19796 11664 19848
rect 11980 19839 12032 19848
rect 11980 19805 11989 19839
rect 11989 19805 12023 19839
rect 12023 19805 12032 19839
rect 11980 19796 12032 19805
rect 12992 19839 13044 19848
rect 12992 19805 13001 19839
rect 13001 19805 13035 19839
rect 13035 19805 13044 19839
rect 15200 19907 15252 19916
rect 15200 19873 15209 19907
rect 15209 19873 15243 19907
rect 15243 19873 15252 19907
rect 15200 19864 15252 19873
rect 15660 19864 15712 19916
rect 12992 19796 13044 19805
rect 16672 19932 16724 19984
rect 24860 19932 24912 19984
rect 11428 19771 11480 19780
rect 11428 19737 11437 19771
rect 11437 19737 11471 19771
rect 11471 19737 11480 19771
rect 11428 19728 11480 19737
rect 9404 19703 9456 19712
rect 9404 19669 9413 19703
rect 9413 19669 9447 19703
rect 9447 19669 9456 19703
rect 9404 19660 9456 19669
rect 10876 19660 10928 19712
rect 13820 19771 13872 19780
rect 13820 19737 13829 19771
rect 13829 19737 13863 19771
rect 13863 19737 13872 19771
rect 13820 19728 13872 19737
rect 14188 19728 14240 19780
rect 15476 19728 15528 19780
rect 12256 19660 12308 19712
rect 15752 19660 15804 19712
rect 16580 19728 16632 19780
rect 16764 19660 16816 19712
rect 8214 19558 8266 19610
rect 8278 19558 8330 19610
rect 8342 19558 8394 19610
rect 8406 19558 8458 19610
rect 8470 19558 8522 19610
rect 16214 19558 16266 19610
rect 16278 19558 16330 19610
rect 16342 19558 16394 19610
rect 16406 19558 16458 19610
rect 16470 19558 16522 19610
rect 24214 19558 24266 19610
rect 24278 19558 24330 19610
rect 24342 19558 24394 19610
rect 24406 19558 24458 19610
rect 24470 19558 24522 19610
rect 5356 19499 5408 19508
rect 5356 19465 5365 19499
rect 5365 19465 5399 19499
rect 5399 19465 5408 19499
rect 5356 19456 5408 19465
rect 5448 19456 5500 19508
rect 7012 19499 7064 19508
rect 7012 19465 7021 19499
rect 7021 19465 7055 19499
rect 7055 19465 7064 19499
rect 7012 19456 7064 19465
rect 9404 19456 9456 19508
rect 11244 19499 11296 19508
rect 11244 19465 11253 19499
rect 11253 19465 11287 19499
rect 11287 19465 11296 19499
rect 11244 19456 11296 19465
rect 12256 19499 12308 19508
rect 12256 19465 12265 19499
rect 12265 19465 12299 19499
rect 12299 19465 12308 19499
rect 12256 19456 12308 19465
rect 13820 19456 13872 19508
rect 4712 19388 4764 19440
rect 8760 19388 8812 19440
rect 10048 19388 10100 19440
rect 10784 19431 10836 19440
rect 10784 19397 10801 19431
rect 10801 19397 10836 19431
rect 10784 19388 10836 19397
rect 11612 19388 11664 19440
rect 15476 19388 15528 19440
rect 4804 19320 4856 19372
rect 5816 19363 5868 19372
rect 5816 19329 5825 19363
rect 5825 19329 5859 19363
rect 5859 19329 5868 19363
rect 5816 19320 5868 19329
rect 7104 19320 7156 19372
rect 7472 19363 7524 19372
rect 7472 19329 7481 19363
rect 7481 19329 7515 19363
rect 7515 19329 7524 19363
rect 7472 19320 7524 19329
rect 8576 19320 8628 19372
rect 9036 19363 9088 19372
rect 9036 19329 9045 19363
rect 9045 19329 9079 19363
rect 9079 19329 9088 19363
rect 9036 19320 9088 19329
rect 10416 19320 10468 19372
rect 10876 19363 10928 19372
rect 10876 19329 10885 19363
rect 10885 19329 10919 19363
rect 10919 19329 10928 19363
rect 10876 19320 10928 19329
rect 11060 19363 11112 19372
rect 11060 19329 11069 19363
rect 11069 19329 11103 19363
rect 11103 19329 11112 19363
rect 11060 19320 11112 19329
rect 11520 19320 11572 19372
rect 5540 19252 5592 19304
rect 9128 19252 9180 19304
rect 9956 19295 10008 19304
rect 9956 19261 9965 19295
rect 9965 19261 9999 19295
rect 9999 19261 10008 19295
rect 9956 19252 10008 19261
rect 5172 19184 5224 19236
rect 7288 19159 7340 19168
rect 7288 19125 7297 19159
rect 7297 19125 7331 19159
rect 7331 19125 7340 19159
rect 7288 19116 7340 19125
rect 9496 19184 9548 19236
rect 11244 19252 11296 19304
rect 11428 19252 11480 19304
rect 10876 19184 10928 19236
rect 12072 19363 12124 19372
rect 12072 19329 12081 19363
rect 12081 19329 12115 19363
rect 12115 19329 12124 19363
rect 12072 19320 12124 19329
rect 12716 19320 12768 19372
rect 14188 19363 14240 19372
rect 14188 19329 14197 19363
rect 14197 19329 14231 19363
rect 14231 19329 14240 19363
rect 14188 19320 14240 19329
rect 15016 19320 15068 19372
rect 15384 19252 15436 19304
rect 16028 19252 16080 19304
rect 16580 19456 16632 19508
rect 16764 19431 16816 19440
rect 16764 19397 16773 19431
rect 16773 19397 16807 19431
rect 16807 19397 16816 19431
rect 16764 19388 16816 19397
rect 16396 19252 16448 19304
rect 17592 19252 17644 19304
rect 25596 19252 25648 19304
rect 16764 19184 16816 19236
rect 12532 19116 12584 19168
rect 24952 19116 25004 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 12214 19014 12266 19066
rect 12278 19014 12330 19066
rect 12342 19014 12394 19066
rect 12406 19014 12458 19066
rect 12470 19014 12522 19066
rect 20214 19014 20266 19066
rect 20278 19014 20330 19066
rect 20342 19014 20394 19066
rect 20406 19014 20458 19066
rect 20470 19014 20522 19066
rect 4804 18955 4856 18964
rect 4804 18921 4813 18955
rect 4813 18921 4847 18955
rect 4847 18921 4856 18955
rect 4804 18912 4856 18921
rect 4896 18912 4948 18964
rect 5816 18912 5868 18964
rect 7104 18955 7156 18964
rect 7104 18921 7113 18955
rect 7113 18921 7147 18955
rect 7147 18921 7156 18955
rect 7104 18912 7156 18921
rect 8576 18955 8628 18964
rect 8576 18921 8585 18955
rect 8585 18921 8619 18955
rect 8619 18921 8628 18955
rect 8576 18912 8628 18921
rect 9036 18955 9088 18964
rect 9036 18921 9045 18955
rect 9045 18921 9079 18955
rect 9079 18921 9088 18955
rect 9036 18912 9088 18921
rect 9680 18912 9732 18964
rect 10508 18912 10560 18964
rect 10876 18912 10928 18964
rect 11152 18912 11204 18964
rect 11888 18912 11940 18964
rect 12348 18912 12400 18964
rect 12624 18912 12676 18964
rect 14188 18912 14240 18964
rect 6828 18844 6880 18896
rect 7748 18819 7800 18828
rect 7748 18785 7757 18819
rect 7757 18785 7791 18819
rect 7791 18785 7800 18819
rect 10048 18887 10100 18896
rect 10048 18853 10057 18887
rect 10057 18853 10091 18887
rect 10091 18853 10100 18887
rect 10048 18844 10100 18853
rect 12072 18844 12124 18896
rect 7748 18776 7800 18785
rect 3240 18708 3292 18760
rect 4528 18708 4580 18760
rect 4068 18640 4120 18692
rect 5724 18751 5776 18760
rect 5724 18717 5733 18751
rect 5733 18717 5767 18751
rect 5767 18717 5776 18751
rect 5724 18708 5776 18717
rect 6552 18708 6604 18760
rect 6920 18708 6972 18760
rect 9588 18776 9640 18828
rect 10140 18708 10192 18760
rect 11244 18751 11296 18760
rect 11244 18717 11253 18751
rect 11253 18717 11287 18751
rect 11287 18717 11296 18751
rect 11244 18708 11296 18717
rect 11612 18776 11664 18828
rect 13084 18844 13136 18896
rect 11520 18751 11572 18760
rect 11520 18717 11529 18751
rect 11529 18717 11563 18751
rect 11563 18717 11572 18751
rect 11520 18708 11572 18717
rect 11704 18751 11756 18760
rect 11704 18717 11713 18751
rect 11713 18717 11747 18751
rect 11747 18717 11756 18751
rect 11704 18708 11756 18717
rect 12256 18708 12308 18760
rect 12348 18751 12400 18760
rect 12348 18717 12357 18751
rect 12357 18717 12391 18751
rect 12391 18717 12400 18751
rect 12348 18708 12400 18717
rect 12440 18751 12492 18760
rect 12440 18717 12449 18751
rect 12449 18717 12483 18751
rect 12483 18717 12492 18751
rect 12440 18708 12492 18717
rect 17592 18776 17644 18828
rect 12624 18708 12676 18760
rect 13360 18708 13412 18760
rect 14004 18708 14056 18760
rect 14556 18751 14608 18760
rect 14556 18717 14565 18751
rect 14565 18717 14599 18751
rect 14599 18717 14608 18751
rect 14556 18708 14608 18717
rect 16764 18751 16816 18760
rect 16764 18717 16773 18751
rect 16773 18717 16807 18751
rect 16807 18717 16816 18751
rect 16764 18708 16816 18717
rect 7840 18640 7892 18692
rect 11152 18640 11204 18692
rect 11428 18683 11480 18692
rect 11428 18649 11445 18683
rect 11445 18649 11480 18683
rect 11428 18640 11480 18649
rect 4436 18572 4488 18624
rect 5816 18572 5868 18624
rect 6460 18572 6512 18624
rect 13268 18640 13320 18692
rect 13636 18572 13688 18624
rect 13820 18572 13872 18624
rect 15200 18683 15252 18692
rect 15200 18649 15209 18683
rect 15209 18649 15243 18683
rect 15243 18649 15252 18683
rect 15200 18640 15252 18649
rect 17500 18708 17552 18760
rect 16948 18615 17000 18624
rect 16948 18581 16957 18615
rect 16957 18581 16991 18615
rect 16991 18581 17000 18615
rect 16948 18572 17000 18581
rect 17224 18615 17276 18624
rect 17224 18581 17233 18615
rect 17233 18581 17267 18615
rect 17267 18581 17276 18615
rect 17224 18572 17276 18581
rect 18144 18572 18196 18624
rect 8214 18470 8266 18522
rect 8278 18470 8330 18522
rect 8342 18470 8394 18522
rect 8406 18470 8458 18522
rect 8470 18470 8522 18522
rect 16214 18470 16266 18522
rect 16278 18470 16330 18522
rect 16342 18470 16394 18522
rect 16406 18470 16458 18522
rect 16470 18470 16522 18522
rect 24214 18470 24266 18522
rect 24278 18470 24330 18522
rect 24342 18470 24394 18522
rect 24406 18470 24458 18522
rect 24470 18470 24522 18522
rect 3240 18411 3292 18420
rect 3240 18377 3249 18411
rect 3249 18377 3283 18411
rect 3283 18377 3292 18411
rect 3240 18368 3292 18377
rect 4068 18368 4120 18420
rect 4252 18232 4304 18284
rect 4620 18368 4672 18420
rect 4712 18368 4764 18420
rect 5724 18368 5776 18420
rect 6552 18368 6604 18420
rect 10876 18368 10928 18420
rect 4436 18343 4488 18352
rect 4436 18309 4445 18343
rect 4445 18309 4479 18343
rect 4479 18309 4488 18343
rect 4436 18300 4488 18309
rect 4528 18164 4580 18216
rect 5080 18207 5132 18216
rect 5080 18173 5089 18207
rect 5089 18173 5123 18207
rect 5123 18173 5132 18207
rect 5080 18164 5132 18173
rect 6828 18275 6880 18284
rect 6828 18241 6837 18275
rect 6837 18241 6871 18275
rect 6871 18241 6880 18275
rect 6828 18232 6880 18241
rect 4712 18096 4764 18148
rect 6736 18164 6788 18216
rect 9680 18232 9732 18284
rect 10508 18300 10560 18352
rect 11428 18300 11480 18352
rect 12256 18411 12308 18420
rect 12256 18377 12265 18411
rect 12265 18377 12299 18411
rect 12299 18377 12308 18411
rect 12256 18368 12308 18377
rect 12348 18368 12400 18420
rect 12992 18368 13044 18420
rect 5816 18096 5868 18148
rect 10140 18164 10192 18216
rect 9864 18096 9916 18148
rect 11520 18232 11572 18284
rect 11612 18275 11664 18284
rect 11612 18241 11621 18275
rect 11621 18241 11655 18275
rect 11655 18241 11664 18275
rect 11612 18232 11664 18241
rect 15200 18368 15252 18420
rect 15476 18368 15528 18420
rect 24860 18368 24912 18420
rect 14280 18300 14332 18352
rect 12072 18232 12124 18284
rect 11152 18096 11204 18148
rect 11336 18096 11388 18148
rect 12716 18232 12768 18284
rect 12808 18275 12860 18284
rect 12808 18241 12817 18275
rect 12817 18241 12851 18275
rect 12851 18241 12860 18275
rect 12808 18232 12860 18241
rect 13176 18232 13228 18284
rect 13636 18275 13688 18284
rect 12624 18096 12676 18148
rect 13636 18241 13644 18275
rect 13644 18241 13678 18275
rect 13678 18241 13688 18275
rect 13636 18232 13688 18241
rect 13728 18275 13780 18284
rect 13728 18241 13737 18275
rect 13737 18241 13771 18275
rect 13771 18241 13780 18275
rect 13728 18232 13780 18241
rect 13820 18232 13872 18284
rect 16948 18300 17000 18352
rect 14556 18275 14608 18284
rect 14556 18241 14565 18275
rect 14565 18241 14599 18275
rect 14599 18241 14608 18275
rect 14556 18232 14608 18241
rect 14372 18164 14424 18216
rect 15200 18275 15252 18284
rect 15200 18241 15209 18275
rect 15209 18241 15243 18275
rect 15243 18241 15252 18275
rect 15200 18232 15252 18241
rect 15476 18275 15528 18284
rect 15476 18241 15485 18275
rect 15485 18241 15519 18275
rect 15519 18241 15528 18275
rect 15476 18232 15528 18241
rect 18144 18343 18196 18352
rect 18144 18309 18153 18343
rect 18153 18309 18187 18343
rect 18187 18309 18196 18343
rect 18144 18300 18196 18309
rect 15384 18164 15436 18216
rect 16028 18207 16080 18216
rect 16028 18173 16037 18207
rect 16037 18173 16071 18207
rect 16071 18173 16080 18207
rect 16028 18164 16080 18173
rect 14556 18096 14608 18148
rect 17960 18096 18012 18148
rect 4068 18028 4120 18080
rect 4252 18028 4304 18080
rect 5356 18028 5408 18080
rect 10692 18028 10744 18080
rect 12072 18028 12124 18080
rect 12716 18071 12768 18080
rect 12716 18037 12725 18071
rect 12725 18037 12759 18071
rect 12759 18037 12768 18071
rect 12716 18028 12768 18037
rect 12992 18028 13044 18080
rect 13360 18028 13412 18080
rect 17500 18028 17552 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 12214 17926 12266 17978
rect 12278 17926 12330 17978
rect 12342 17926 12394 17978
rect 12406 17926 12458 17978
rect 12470 17926 12522 17978
rect 20214 17926 20266 17978
rect 20278 17926 20330 17978
rect 20342 17926 20394 17978
rect 20406 17926 20458 17978
rect 20470 17926 20522 17978
rect 4988 17824 5040 17876
rect 5356 17867 5408 17876
rect 5356 17833 5365 17867
rect 5365 17833 5399 17867
rect 5399 17833 5408 17867
rect 5356 17824 5408 17833
rect 4344 17756 4396 17808
rect 5080 17756 5132 17808
rect 10324 17824 10376 17876
rect 4436 17663 4488 17672
rect 4436 17629 4445 17663
rect 4445 17629 4479 17663
rect 4479 17629 4488 17663
rect 4436 17620 4488 17629
rect 7288 17688 7340 17740
rect 4712 17620 4764 17672
rect 4344 17552 4396 17604
rect 5632 17663 5684 17672
rect 5632 17629 5641 17663
rect 5641 17629 5675 17663
rect 5675 17629 5684 17663
rect 5632 17620 5684 17629
rect 5816 17620 5868 17672
rect 6552 17620 6604 17672
rect 7012 17620 7064 17672
rect 8576 17620 8628 17672
rect 9404 17756 9456 17808
rect 11428 17824 11480 17876
rect 11520 17867 11572 17876
rect 11520 17833 11529 17867
rect 11529 17833 11563 17867
rect 11563 17833 11572 17867
rect 11520 17824 11572 17833
rect 11888 17824 11940 17876
rect 10232 17688 10284 17740
rect 9772 17620 9824 17672
rect 10600 17756 10652 17808
rect 12992 17824 13044 17876
rect 13084 17824 13136 17876
rect 12716 17756 12768 17808
rect 12808 17756 12860 17808
rect 13268 17756 13320 17808
rect 15568 17824 15620 17876
rect 16028 17824 16080 17876
rect 15476 17756 15528 17808
rect 17224 17756 17276 17808
rect 10416 17663 10468 17672
rect 10416 17629 10425 17663
rect 10425 17629 10459 17663
rect 10459 17629 10468 17663
rect 10416 17620 10468 17629
rect 10600 17663 10652 17672
rect 10600 17629 10609 17663
rect 10609 17629 10643 17663
rect 10643 17629 10652 17663
rect 10600 17620 10652 17629
rect 10968 17620 11020 17672
rect 10140 17595 10192 17604
rect 10140 17561 10149 17595
rect 10149 17561 10183 17595
rect 10183 17561 10192 17595
rect 10140 17552 10192 17561
rect 4436 17484 4488 17536
rect 5816 17484 5868 17536
rect 6184 17484 6236 17536
rect 7564 17527 7616 17536
rect 7564 17493 7573 17527
rect 7573 17493 7607 17527
rect 7607 17493 7616 17527
rect 7564 17484 7616 17493
rect 7932 17484 7984 17536
rect 10784 17552 10836 17604
rect 11152 17552 11204 17604
rect 12716 17620 12768 17672
rect 13820 17688 13872 17740
rect 12992 17663 13044 17672
rect 12992 17629 13001 17663
rect 13001 17629 13035 17663
rect 13035 17629 13044 17663
rect 12992 17620 13044 17629
rect 13452 17663 13504 17672
rect 13452 17629 13461 17663
rect 13461 17629 13495 17663
rect 13495 17629 13504 17663
rect 13452 17620 13504 17629
rect 13636 17620 13688 17672
rect 10876 17527 10928 17536
rect 10876 17493 10885 17527
rect 10885 17493 10919 17527
rect 10919 17493 10928 17527
rect 10876 17484 10928 17493
rect 11796 17484 11848 17536
rect 12164 17527 12216 17536
rect 12164 17493 12173 17527
rect 12173 17493 12207 17527
rect 12207 17493 12216 17527
rect 12164 17484 12216 17493
rect 12256 17484 12308 17536
rect 12808 17484 12860 17536
rect 12900 17527 12952 17536
rect 12900 17493 12909 17527
rect 12909 17493 12943 17527
rect 12943 17493 12952 17527
rect 12900 17484 12952 17493
rect 12992 17484 13044 17536
rect 13820 17552 13872 17604
rect 14372 17620 14424 17672
rect 14648 17663 14700 17672
rect 14648 17629 14662 17663
rect 14662 17629 14696 17663
rect 14696 17629 14700 17663
rect 14648 17620 14700 17629
rect 15568 17663 15620 17672
rect 15568 17629 15577 17663
rect 15577 17629 15611 17663
rect 15611 17629 15620 17663
rect 15568 17620 15620 17629
rect 16028 17620 16080 17672
rect 14464 17595 14516 17604
rect 14464 17561 14473 17595
rect 14473 17561 14507 17595
rect 14507 17561 14516 17595
rect 14464 17552 14516 17561
rect 13912 17484 13964 17536
rect 14280 17484 14332 17536
rect 15936 17552 15988 17604
rect 17960 17663 18012 17672
rect 17960 17629 17969 17663
rect 17969 17629 18003 17663
rect 18003 17629 18012 17663
rect 17960 17620 18012 17629
rect 18236 17552 18288 17604
rect 14832 17527 14884 17536
rect 14832 17493 14841 17527
rect 14841 17493 14875 17527
rect 14875 17493 14884 17527
rect 14832 17484 14884 17493
rect 16120 17484 16172 17536
rect 17500 17484 17552 17536
rect 18420 17527 18472 17536
rect 18420 17493 18429 17527
rect 18429 17493 18463 17527
rect 18463 17493 18472 17527
rect 18420 17484 18472 17493
rect 8214 17382 8266 17434
rect 8278 17382 8330 17434
rect 8342 17382 8394 17434
rect 8406 17382 8458 17434
rect 8470 17382 8522 17434
rect 16214 17382 16266 17434
rect 16278 17382 16330 17434
rect 16342 17382 16394 17434
rect 16406 17382 16458 17434
rect 16470 17382 16522 17434
rect 24214 17382 24266 17434
rect 24278 17382 24330 17434
rect 24342 17382 24394 17434
rect 24406 17382 24458 17434
rect 24470 17382 24522 17434
rect 4712 17323 4764 17332
rect 4712 17289 4721 17323
rect 4721 17289 4755 17323
rect 4755 17289 4764 17323
rect 4712 17280 4764 17289
rect 4344 17255 4396 17264
rect 4344 17221 4353 17255
rect 4353 17221 4387 17255
rect 4387 17221 4396 17255
rect 4344 17212 4396 17221
rect 4436 17255 4488 17264
rect 4436 17221 4445 17255
rect 4445 17221 4479 17255
rect 4479 17221 4488 17255
rect 4436 17212 4488 17221
rect 4528 17212 4580 17264
rect 4988 17144 5040 17196
rect 7012 17255 7064 17264
rect 7012 17221 7021 17255
rect 7021 17221 7055 17255
rect 7055 17221 7064 17255
rect 7012 17212 7064 17221
rect 5816 17144 5868 17196
rect 6092 17144 6144 17196
rect 7564 17144 7616 17196
rect 7932 17187 7984 17196
rect 7932 17153 7941 17187
rect 7941 17153 7975 17187
rect 7975 17153 7984 17187
rect 7932 17144 7984 17153
rect 8392 17187 8444 17196
rect 8392 17153 8401 17187
rect 8401 17153 8435 17187
rect 8435 17153 8444 17187
rect 8392 17144 8444 17153
rect 3884 17119 3936 17128
rect 3884 17085 3893 17119
rect 3893 17085 3927 17119
rect 3927 17085 3936 17119
rect 3884 17076 3936 17085
rect 4712 17119 4764 17128
rect 4712 17085 4721 17119
rect 4721 17085 4755 17119
rect 4755 17085 4764 17119
rect 4712 17076 4764 17085
rect 7472 17119 7524 17128
rect 7472 17085 7481 17119
rect 7481 17085 7515 17119
rect 7515 17085 7524 17119
rect 7472 17076 7524 17085
rect 8484 17076 8536 17128
rect 5908 16983 5960 16992
rect 5908 16949 5917 16983
rect 5917 16949 5951 16983
rect 5951 16949 5960 16983
rect 5908 16940 5960 16949
rect 7840 16940 7892 16992
rect 9128 17187 9180 17196
rect 9128 17153 9137 17187
rect 9137 17153 9171 17187
rect 9171 17153 9180 17187
rect 9128 17144 9180 17153
rect 10876 17280 10928 17332
rect 12164 17280 12216 17332
rect 12900 17280 12952 17332
rect 14004 17280 14056 17332
rect 14096 17280 14148 17332
rect 9404 17187 9456 17196
rect 9404 17153 9413 17187
rect 9413 17153 9447 17187
rect 9447 17153 9456 17187
rect 9404 17144 9456 17153
rect 9680 17187 9732 17196
rect 9680 17153 9689 17187
rect 9689 17153 9723 17187
rect 9723 17153 9732 17187
rect 9680 17144 9732 17153
rect 9864 17187 9916 17196
rect 9864 17153 9873 17187
rect 9873 17153 9907 17187
rect 9907 17153 9916 17187
rect 9864 17144 9916 17153
rect 9956 17187 10008 17196
rect 9956 17153 9965 17187
rect 9965 17153 9999 17187
rect 9999 17153 10008 17187
rect 9956 17144 10008 17153
rect 10140 17144 10192 17196
rect 10508 17144 10560 17196
rect 10600 17187 10652 17196
rect 10600 17153 10609 17187
rect 10609 17153 10643 17187
rect 10643 17153 10652 17187
rect 10600 17144 10652 17153
rect 11244 17144 11296 17196
rect 11428 17144 11480 17196
rect 12624 17144 12676 17196
rect 12808 17187 12860 17196
rect 12808 17153 12817 17187
rect 12817 17153 12851 17187
rect 12851 17153 12860 17187
rect 12808 17144 12860 17153
rect 12900 17187 12952 17196
rect 12900 17153 12909 17187
rect 12909 17153 12943 17187
rect 12943 17153 12952 17187
rect 12900 17144 12952 17153
rect 9128 17008 9180 17060
rect 9496 17008 9548 17060
rect 9956 17008 10008 17060
rect 10048 16940 10100 16992
rect 10232 17051 10284 17060
rect 10232 17017 10241 17051
rect 10241 17017 10275 17051
rect 10275 17017 10284 17051
rect 10232 17008 10284 17017
rect 10968 17008 11020 17060
rect 11336 17008 11388 17060
rect 11612 17051 11664 17060
rect 11612 17017 11621 17051
rect 11621 17017 11655 17051
rect 11655 17017 11664 17051
rect 11612 17008 11664 17017
rect 12072 17076 12124 17128
rect 13268 17119 13320 17128
rect 13268 17085 13277 17119
rect 13277 17085 13311 17119
rect 13311 17085 13320 17119
rect 13268 17076 13320 17085
rect 13452 17187 13504 17196
rect 13452 17153 13461 17187
rect 13461 17153 13495 17187
rect 13495 17153 13504 17187
rect 13452 17144 13504 17153
rect 13728 17144 13780 17196
rect 14280 17255 14332 17264
rect 14280 17221 14289 17255
rect 14289 17221 14323 17255
rect 14323 17221 14332 17255
rect 14280 17212 14332 17221
rect 14188 17187 14240 17196
rect 14188 17153 14197 17187
rect 14197 17153 14231 17187
rect 14231 17153 14240 17187
rect 14188 17144 14240 17153
rect 14832 17212 14884 17264
rect 16948 17187 17000 17196
rect 16948 17153 16956 17187
rect 16956 17153 17000 17187
rect 16948 17144 17000 17153
rect 18236 17187 18288 17196
rect 18236 17153 18245 17187
rect 18245 17153 18279 17187
rect 18279 17153 18288 17187
rect 18236 17144 18288 17153
rect 19340 17187 19392 17196
rect 19340 17153 19349 17187
rect 19349 17153 19383 17187
rect 19383 17153 19392 17187
rect 19340 17144 19392 17153
rect 11980 17008 12032 17060
rect 12164 17008 12216 17060
rect 17132 17008 17184 17060
rect 19524 17008 19576 17060
rect 14556 16983 14608 16992
rect 14556 16949 14565 16983
rect 14565 16949 14599 16983
rect 14599 16949 14608 16983
rect 14556 16940 14608 16949
rect 16580 16940 16632 16992
rect 17040 16940 17092 16992
rect 21548 16940 21600 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 12214 16838 12266 16890
rect 12278 16838 12330 16890
rect 12342 16838 12394 16890
rect 12406 16838 12458 16890
rect 12470 16838 12522 16890
rect 20214 16838 20266 16890
rect 20278 16838 20330 16890
rect 20342 16838 20394 16890
rect 20406 16838 20458 16890
rect 20470 16838 20522 16890
rect 3884 16736 3936 16788
rect 4712 16736 4764 16788
rect 7012 16736 7064 16788
rect 8576 16736 8628 16788
rect 11520 16736 11572 16788
rect 11612 16779 11664 16788
rect 11612 16745 11621 16779
rect 11621 16745 11655 16779
rect 11655 16745 11664 16779
rect 11612 16736 11664 16745
rect 11888 16736 11940 16788
rect 23572 16736 23624 16788
rect 3976 16575 4028 16584
rect 3976 16541 3985 16575
rect 3985 16541 4019 16575
rect 4019 16541 4028 16575
rect 3976 16532 4028 16541
rect 4252 16575 4304 16584
rect 4252 16541 4261 16575
rect 4261 16541 4295 16575
rect 4295 16541 4304 16575
rect 4252 16532 4304 16541
rect 4988 16575 5040 16584
rect 4988 16541 4997 16575
rect 4997 16541 5031 16575
rect 5031 16541 5040 16575
rect 5908 16668 5960 16720
rect 4988 16532 5040 16541
rect 5816 16532 5868 16584
rect 7472 16600 7524 16652
rect 7288 16532 7340 16584
rect 7380 16575 7432 16584
rect 7380 16541 7389 16575
rect 7389 16541 7423 16575
rect 7423 16541 7432 16575
rect 7380 16532 7432 16541
rect 7656 16575 7708 16584
rect 7656 16541 7665 16575
rect 7665 16541 7699 16575
rect 7699 16541 7708 16575
rect 7656 16532 7708 16541
rect 8392 16532 8444 16584
rect 6276 16507 6328 16516
rect 6276 16473 6285 16507
rect 6285 16473 6319 16507
rect 6319 16473 6328 16507
rect 6276 16464 6328 16473
rect 7748 16464 7800 16516
rect 8760 16532 8812 16584
rect 9312 16600 9364 16652
rect 9588 16600 9640 16652
rect 11980 16668 12032 16720
rect 12256 16668 12308 16720
rect 8852 16464 8904 16516
rect 9128 16464 9180 16516
rect 4160 16396 4212 16448
rect 5724 16396 5776 16448
rect 9680 16464 9732 16516
rect 10140 16575 10192 16584
rect 10140 16541 10149 16575
rect 10149 16541 10183 16575
rect 10183 16541 10192 16575
rect 10140 16532 10192 16541
rect 10508 16575 10560 16584
rect 10508 16541 10517 16575
rect 10517 16541 10551 16575
rect 10551 16541 10560 16575
rect 10508 16532 10560 16541
rect 10876 16532 10928 16584
rect 11612 16600 11664 16652
rect 12624 16668 12676 16720
rect 12808 16668 12860 16720
rect 12992 16668 13044 16720
rect 14924 16668 14976 16720
rect 16028 16668 16080 16720
rect 11336 16575 11388 16584
rect 11336 16541 11345 16575
rect 11345 16541 11379 16575
rect 11379 16541 11388 16575
rect 11336 16532 11388 16541
rect 11520 16532 11572 16584
rect 12164 16575 12216 16584
rect 12164 16541 12173 16575
rect 12173 16541 12207 16575
rect 12207 16541 12216 16575
rect 12164 16532 12216 16541
rect 12532 16532 12584 16584
rect 12808 16575 12860 16584
rect 12808 16541 12817 16575
rect 12817 16541 12851 16575
rect 12851 16541 12860 16575
rect 12808 16532 12860 16541
rect 13544 16600 13596 16652
rect 13176 16532 13228 16584
rect 13728 16532 13780 16584
rect 15108 16575 15160 16584
rect 15108 16541 15117 16575
rect 15117 16541 15151 16575
rect 15151 16541 15160 16575
rect 15108 16532 15160 16541
rect 15752 16532 15804 16584
rect 16764 16643 16816 16652
rect 16764 16609 16773 16643
rect 16773 16609 16807 16643
rect 16807 16609 16816 16643
rect 16764 16600 16816 16609
rect 16948 16711 17000 16720
rect 16948 16677 16957 16711
rect 16957 16677 16991 16711
rect 16991 16677 17000 16711
rect 16948 16668 17000 16677
rect 18420 16711 18472 16720
rect 18420 16677 18429 16711
rect 18429 16677 18463 16711
rect 18463 16677 18472 16711
rect 18420 16668 18472 16677
rect 16212 16575 16264 16584
rect 16212 16541 16221 16575
rect 16221 16541 16255 16575
rect 16255 16541 16264 16575
rect 16212 16532 16264 16541
rect 12072 16464 12124 16516
rect 12256 16464 12308 16516
rect 15384 16464 15436 16516
rect 17132 16507 17184 16516
rect 17132 16473 17141 16507
rect 17141 16473 17175 16507
rect 17175 16473 17184 16507
rect 17132 16464 17184 16473
rect 18236 16532 18288 16584
rect 19340 16532 19392 16584
rect 26148 16464 26200 16516
rect 9496 16396 9548 16448
rect 11244 16396 11296 16448
rect 11796 16396 11848 16448
rect 12440 16439 12492 16448
rect 12440 16405 12449 16439
rect 12449 16405 12483 16439
rect 12483 16405 12492 16439
rect 12440 16396 12492 16405
rect 16764 16396 16816 16448
rect 8214 16294 8266 16346
rect 8278 16294 8330 16346
rect 8342 16294 8394 16346
rect 8406 16294 8458 16346
rect 8470 16294 8522 16346
rect 16214 16294 16266 16346
rect 16278 16294 16330 16346
rect 16342 16294 16394 16346
rect 16406 16294 16458 16346
rect 16470 16294 16522 16346
rect 24214 16294 24266 16346
rect 24278 16294 24330 16346
rect 24342 16294 24394 16346
rect 24406 16294 24458 16346
rect 24470 16294 24522 16346
rect 7656 16192 7708 16244
rect 8852 16192 8904 16244
rect 9496 16192 9548 16244
rect 10784 16192 10836 16244
rect 11612 16235 11664 16244
rect 11612 16201 11621 16235
rect 11621 16201 11655 16235
rect 11655 16201 11664 16235
rect 11612 16192 11664 16201
rect 11796 16192 11848 16244
rect 12992 16192 13044 16244
rect 13268 16192 13320 16244
rect 13360 16235 13412 16244
rect 13360 16201 13369 16235
rect 13369 16201 13403 16235
rect 13403 16201 13412 16235
rect 13360 16192 13412 16201
rect 14188 16235 14240 16244
rect 14188 16201 14197 16235
rect 14197 16201 14231 16235
rect 14231 16201 14240 16235
rect 14188 16192 14240 16201
rect 15108 16192 15160 16244
rect 4252 16124 4304 16176
rect 10508 16124 10560 16176
rect 11980 16124 12032 16176
rect 12532 16124 12584 16176
rect 3056 15988 3108 16040
rect 3424 16099 3476 16108
rect 3424 16065 3433 16099
rect 3433 16065 3467 16099
rect 3467 16065 3476 16099
rect 4160 16099 4212 16108
rect 3424 16056 3476 16065
rect 4160 16065 4169 16099
rect 4169 16065 4203 16099
rect 4203 16065 4212 16099
rect 4160 16056 4212 16065
rect 6092 16099 6144 16108
rect 6092 16065 6101 16099
rect 6101 16065 6135 16099
rect 6135 16065 6144 16099
rect 6092 16056 6144 16065
rect 8300 16056 8352 16108
rect 9128 16056 9180 16108
rect 9220 16099 9272 16108
rect 9220 16065 9229 16099
rect 9229 16065 9263 16099
rect 9263 16065 9272 16099
rect 9220 16056 9272 16065
rect 9312 16056 9364 16108
rect 10692 16056 10744 16108
rect 10232 15988 10284 16040
rect 3148 15852 3200 15904
rect 4620 15852 4672 15904
rect 6092 15895 6144 15904
rect 6092 15861 6101 15895
rect 6101 15861 6135 15895
rect 6135 15861 6144 15895
rect 6092 15852 6144 15861
rect 7748 15920 7800 15972
rect 9588 15920 9640 15972
rect 10048 15963 10100 15972
rect 10048 15929 10057 15963
rect 10057 15929 10091 15963
rect 10091 15929 10100 15963
rect 10048 15920 10100 15929
rect 11336 16056 11388 16108
rect 11428 16056 11480 16108
rect 11152 15988 11204 16040
rect 12440 16056 12492 16108
rect 12716 16099 12768 16108
rect 12716 16065 12725 16099
rect 12725 16065 12759 16099
rect 12759 16065 12768 16099
rect 12716 16056 12768 16065
rect 12808 16099 12860 16108
rect 12808 16065 12817 16099
rect 12817 16065 12851 16099
rect 12851 16065 12860 16099
rect 14556 16124 14608 16176
rect 15568 16124 15620 16176
rect 16212 16124 16264 16176
rect 12808 16056 12860 16065
rect 15108 16056 15160 16108
rect 12072 16031 12124 16040
rect 12072 15997 12081 16031
rect 12081 15997 12115 16031
rect 12115 15997 12124 16031
rect 12072 15988 12124 15997
rect 12900 16031 12952 16040
rect 11520 15920 11572 15972
rect 12900 15997 12909 16031
rect 12909 15997 12943 16031
rect 12943 15997 12952 16031
rect 12900 15988 12952 15997
rect 13728 15988 13780 16040
rect 16948 16192 17000 16244
rect 16764 16099 16816 16108
rect 16764 16065 16773 16099
rect 16773 16065 16807 16099
rect 16807 16065 16816 16099
rect 16764 16056 16816 16065
rect 17132 16056 17184 16108
rect 26424 15988 26476 16040
rect 8024 15852 8076 15904
rect 9864 15852 9916 15904
rect 10324 15852 10376 15904
rect 11704 15852 11756 15904
rect 12992 15852 13044 15904
rect 17316 15852 17368 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 12214 15750 12266 15802
rect 12278 15750 12330 15802
rect 12342 15750 12394 15802
rect 12406 15750 12458 15802
rect 12470 15750 12522 15802
rect 20214 15750 20266 15802
rect 20278 15750 20330 15802
rect 20342 15750 20394 15802
rect 20406 15750 20458 15802
rect 20470 15750 20522 15802
rect 3424 15648 3476 15700
rect 6276 15648 6328 15700
rect 3056 15580 3108 15632
rect 5724 15580 5776 15632
rect 9220 15648 9272 15700
rect 3240 15555 3292 15564
rect 3240 15521 3249 15555
rect 3249 15521 3283 15555
rect 3283 15521 3292 15555
rect 3240 15512 3292 15521
rect 3056 15444 3108 15496
rect 3884 15487 3936 15496
rect 3884 15453 3893 15487
rect 3893 15453 3927 15487
rect 3927 15453 3936 15487
rect 3884 15444 3936 15453
rect 6092 15444 6144 15496
rect 8024 15487 8076 15496
rect 8024 15453 8033 15487
rect 8033 15453 8067 15487
rect 8067 15453 8076 15487
rect 8024 15444 8076 15453
rect 8668 15512 8720 15564
rect 9772 15580 9824 15632
rect 10416 15580 10468 15632
rect 11060 15648 11112 15700
rect 12900 15648 12952 15700
rect 10968 15580 11020 15632
rect 8576 15444 8628 15496
rect 9404 15444 9456 15496
rect 10232 15512 10284 15564
rect 12440 15580 12492 15632
rect 13084 15580 13136 15632
rect 11336 15512 11388 15564
rect 13728 15512 13780 15564
rect 14556 15512 14608 15564
rect 16212 15555 16264 15564
rect 16212 15521 16221 15555
rect 16221 15521 16255 15555
rect 16255 15521 16264 15555
rect 16212 15512 16264 15521
rect 2964 15308 3016 15360
rect 4620 15376 4672 15428
rect 8300 15376 8352 15428
rect 8852 15376 8904 15428
rect 9588 15376 9640 15428
rect 4988 15308 5040 15360
rect 8116 15351 8168 15360
rect 8116 15317 8125 15351
rect 8125 15317 8159 15351
rect 8159 15317 8168 15351
rect 8116 15308 8168 15317
rect 10324 15376 10376 15428
rect 11244 15444 11296 15496
rect 11704 15487 11756 15496
rect 11704 15453 11713 15487
rect 11713 15453 11747 15487
rect 11747 15453 11756 15487
rect 11704 15444 11756 15453
rect 11888 15487 11940 15496
rect 11888 15453 11897 15487
rect 11897 15453 11931 15487
rect 11931 15453 11940 15487
rect 11888 15444 11940 15453
rect 12716 15444 12768 15496
rect 13636 15487 13688 15496
rect 13636 15453 13645 15487
rect 13645 15453 13679 15487
rect 13679 15453 13688 15487
rect 13636 15444 13688 15453
rect 16580 15444 16632 15496
rect 10140 15308 10192 15360
rect 11152 15351 11204 15360
rect 11152 15317 11161 15351
rect 11161 15317 11195 15351
rect 11195 15317 11204 15351
rect 11152 15308 11204 15317
rect 13084 15376 13136 15428
rect 13176 15419 13228 15428
rect 13176 15385 13185 15419
rect 13185 15385 13219 15419
rect 13219 15385 13228 15419
rect 13176 15376 13228 15385
rect 12808 15308 12860 15360
rect 8214 15206 8266 15258
rect 8278 15206 8330 15258
rect 8342 15206 8394 15258
rect 8406 15206 8458 15258
rect 8470 15206 8522 15258
rect 16214 15206 16266 15258
rect 16278 15206 16330 15258
rect 16342 15206 16394 15258
rect 16406 15206 16458 15258
rect 16470 15206 16522 15258
rect 24214 15206 24266 15258
rect 24278 15206 24330 15258
rect 24342 15206 24394 15258
rect 24406 15206 24458 15258
rect 24470 15206 24522 15258
rect 1492 14900 1544 14952
rect 3884 15104 3936 15156
rect 6828 15104 6880 15156
rect 2964 15036 3016 15088
rect 3240 15036 3292 15088
rect 4068 15036 4120 15088
rect 8116 15036 8168 15088
rect 8576 15147 8628 15156
rect 8576 15113 8585 15147
rect 8585 15113 8619 15147
rect 8619 15113 8628 15147
rect 8576 15104 8628 15113
rect 10048 15147 10100 15156
rect 10048 15113 10057 15147
rect 10057 15113 10091 15147
rect 10091 15113 10100 15147
rect 10048 15104 10100 15113
rect 10876 15104 10928 15156
rect 11428 15104 11480 15156
rect 11980 15104 12032 15156
rect 12808 15147 12860 15156
rect 12808 15113 12817 15147
rect 12817 15113 12851 15147
rect 12851 15113 12860 15147
rect 12808 15104 12860 15113
rect 9864 15036 9916 15088
rect 3976 14968 4028 15020
rect 4804 14968 4856 15020
rect 2688 14900 2740 14952
rect 3240 14900 3292 14952
rect 5080 14943 5132 14952
rect 5080 14909 5089 14943
rect 5089 14909 5123 14943
rect 5123 14909 5132 14943
rect 5080 14900 5132 14909
rect 9128 14968 9180 15020
rect 10048 15011 10100 15020
rect 10048 14977 10057 15011
rect 10057 14977 10091 15011
rect 10091 14977 10100 15011
rect 10048 14968 10100 14977
rect 10232 15011 10284 15020
rect 10232 14977 10241 15011
rect 10241 14977 10275 15011
rect 10275 14977 10284 15011
rect 10232 14968 10284 14977
rect 11152 14968 11204 15020
rect 11244 15011 11296 15020
rect 11244 14977 11253 15011
rect 11253 14977 11287 15011
rect 11287 14977 11296 15011
rect 11244 14968 11296 14977
rect 11336 14968 11388 15020
rect 12072 14968 12124 15020
rect 13176 15036 13228 15088
rect 16120 15079 16172 15088
rect 16120 15045 16129 15079
rect 16129 15045 16163 15079
rect 16163 15045 16172 15079
rect 16120 15036 16172 15045
rect 4988 14832 5040 14884
rect 3424 14807 3476 14816
rect 3424 14773 3433 14807
rect 3433 14773 3467 14807
rect 3467 14773 3476 14807
rect 3424 14764 3476 14773
rect 3516 14764 3568 14816
rect 5724 14764 5776 14816
rect 6828 14943 6880 14952
rect 6828 14909 6837 14943
rect 6837 14909 6871 14943
rect 6871 14909 6880 14943
rect 6828 14900 6880 14909
rect 7104 14943 7156 14952
rect 7104 14909 7113 14943
rect 7113 14909 7147 14943
rect 7147 14909 7156 14943
rect 7104 14900 7156 14909
rect 9680 14900 9732 14952
rect 13728 15011 13780 15020
rect 13728 14977 13737 15011
rect 13737 14977 13771 15011
rect 13771 14977 13780 15011
rect 13728 14968 13780 14977
rect 16304 15011 16356 15020
rect 16304 14977 16313 15011
rect 16313 14977 16347 15011
rect 16347 14977 16356 15011
rect 16304 14968 16356 14977
rect 16948 15011 17000 15020
rect 16948 14977 16957 15011
rect 16957 14977 16991 15011
rect 16991 14977 17000 15011
rect 16948 14968 17000 14977
rect 15108 14900 15160 14952
rect 9312 14832 9364 14884
rect 7840 14764 7892 14816
rect 12716 14832 12768 14884
rect 13636 14832 13688 14884
rect 12624 14764 12676 14816
rect 16856 14807 16908 14816
rect 16856 14773 16865 14807
rect 16865 14773 16899 14807
rect 16899 14773 16908 14807
rect 16856 14764 16908 14773
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 12214 14662 12266 14714
rect 12278 14662 12330 14714
rect 12342 14662 12394 14714
rect 12406 14662 12458 14714
rect 12470 14662 12522 14714
rect 20214 14662 20266 14714
rect 20278 14662 20330 14714
rect 20342 14662 20394 14714
rect 20406 14662 20458 14714
rect 20470 14662 20522 14714
rect 4068 14560 4120 14612
rect 3056 14492 3108 14544
rect 2136 14424 2188 14476
rect 1492 14356 1544 14408
rect 3148 14356 3200 14408
rect 4068 14399 4120 14408
rect 4068 14365 4077 14399
rect 4077 14365 4111 14399
rect 4111 14365 4120 14399
rect 4068 14356 4120 14365
rect 5080 14603 5132 14612
rect 5080 14569 5089 14603
rect 5089 14569 5123 14603
rect 5123 14569 5132 14603
rect 5080 14560 5132 14569
rect 7104 14560 7156 14612
rect 8668 14560 8720 14612
rect 9680 14560 9732 14612
rect 9864 14560 9916 14612
rect 2964 14220 3016 14272
rect 3608 14220 3660 14272
rect 3884 14263 3936 14272
rect 3884 14229 3893 14263
rect 3893 14229 3927 14263
rect 3927 14229 3936 14263
rect 3884 14220 3936 14229
rect 4988 14356 5040 14408
rect 5264 14288 5316 14340
rect 5356 14288 5408 14340
rect 6092 14399 6144 14408
rect 6092 14365 6101 14399
rect 6101 14365 6135 14399
rect 6135 14365 6144 14399
rect 6092 14356 6144 14365
rect 6644 14399 6696 14408
rect 6644 14365 6653 14399
rect 6653 14365 6687 14399
rect 6687 14365 6696 14399
rect 6644 14356 6696 14365
rect 8576 14424 8628 14476
rect 9312 14467 9364 14476
rect 9312 14433 9321 14467
rect 9321 14433 9355 14467
rect 9355 14433 9364 14467
rect 9312 14424 9364 14433
rect 11060 14492 11112 14544
rect 9772 14467 9824 14476
rect 9772 14433 9781 14467
rect 9781 14433 9815 14467
rect 9815 14433 9824 14467
rect 9772 14424 9824 14433
rect 7288 14399 7340 14408
rect 7288 14365 7297 14399
rect 7297 14365 7331 14399
rect 7331 14365 7340 14399
rect 7288 14356 7340 14365
rect 6828 14288 6880 14340
rect 8852 14356 8904 14408
rect 9220 14356 9272 14408
rect 10324 14356 10376 14408
rect 10784 14424 10836 14476
rect 11888 14492 11940 14544
rect 12624 14560 12676 14612
rect 13728 14560 13780 14612
rect 15752 14560 15804 14612
rect 16948 14560 17000 14612
rect 8944 14288 8996 14340
rect 9036 14288 9088 14340
rect 10784 14288 10836 14340
rect 12716 14399 12768 14408
rect 12716 14365 12725 14399
rect 12725 14365 12759 14399
rect 12759 14365 12768 14399
rect 12716 14356 12768 14365
rect 12808 14399 12860 14408
rect 12808 14365 12817 14399
rect 12817 14365 12851 14399
rect 12851 14365 12860 14399
rect 12808 14356 12860 14365
rect 12900 14399 12952 14408
rect 12900 14365 12909 14399
rect 12909 14365 12943 14399
rect 12943 14365 12952 14399
rect 12900 14356 12952 14365
rect 14464 14424 14516 14476
rect 16304 14467 16356 14476
rect 16304 14433 16313 14467
rect 16313 14433 16347 14467
rect 16347 14433 16356 14467
rect 16304 14424 16356 14433
rect 13268 14356 13320 14408
rect 14188 14399 14240 14408
rect 14188 14365 14197 14399
rect 14197 14365 14231 14399
rect 14231 14365 14240 14399
rect 14188 14356 14240 14365
rect 15752 14356 15804 14408
rect 15844 14399 15896 14408
rect 15844 14365 15853 14399
rect 15853 14365 15887 14399
rect 15887 14365 15896 14399
rect 15844 14356 15896 14365
rect 16120 14356 16172 14408
rect 12624 14288 12676 14340
rect 13084 14288 13136 14340
rect 13176 14288 13228 14340
rect 4988 14220 5040 14272
rect 5816 14220 5868 14272
rect 7748 14263 7800 14272
rect 7748 14229 7757 14263
rect 7757 14229 7791 14263
rect 7791 14229 7800 14263
rect 7748 14220 7800 14229
rect 9128 14263 9180 14272
rect 9128 14229 9137 14263
rect 9137 14229 9171 14263
rect 9171 14229 9180 14263
rect 9128 14220 9180 14229
rect 11060 14220 11112 14272
rect 11244 14220 11296 14272
rect 11980 14263 12032 14272
rect 11980 14229 11989 14263
rect 11989 14229 12023 14263
rect 12023 14229 12032 14263
rect 11980 14220 12032 14229
rect 14372 14263 14424 14272
rect 14372 14229 14381 14263
rect 14381 14229 14415 14263
rect 14415 14229 14424 14263
rect 14372 14220 14424 14229
rect 8214 14118 8266 14170
rect 8278 14118 8330 14170
rect 8342 14118 8394 14170
rect 8406 14118 8458 14170
rect 8470 14118 8522 14170
rect 16214 14118 16266 14170
rect 16278 14118 16330 14170
rect 16342 14118 16394 14170
rect 16406 14118 16458 14170
rect 16470 14118 16522 14170
rect 24214 14118 24266 14170
rect 24278 14118 24330 14170
rect 24342 14118 24394 14170
rect 24406 14118 24458 14170
rect 24470 14118 24522 14170
rect 3056 14016 3108 14068
rect 3884 14016 3936 14068
rect 3516 13948 3568 14000
rect 3608 13948 3660 14000
rect 5264 14016 5316 14068
rect 6644 14016 6696 14068
rect 7748 14016 7800 14068
rect 4068 13948 4120 14000
rect 2136 13923 2188 13932
rect 2136 13889 2145 13923
rect 2145 13889 2179 13923
rect 2179 13889 2188 13923
rect 2136 13880 2188 13889
rect 4160 13880 4212 13932
rect 2688 13855 2740 13864
rect 2688 13821 2697 13855
rect 2697 13821 2731 13855
rect 2731 13821 2740 13855
rect 2688 13812 2740 13821
rect 3424 13812 3476 13864
rect 3332 13744 3384 13796
rect 4620 13812 4672 13864
rect 4804 13855 4856 13864
rect 4804 13821 4813 13855
rect 4813 13821 4847 13855
rect 4847 13821 4856 13855
rect 4804 13812 4856 13821
rect 6092 13948 6144 14000
rect 6828 13991 6880 14000
rect 6828 13957 6837 13991
rect 6837 13957 6871 13991
rect 6871 13957 6880 13991
rect 6828 13948 6880 13957
rect 5264 13880 5316 13932
rect 5724 13923 5776 13932
rect 5724 13889 5733 13923
rect 5733 13889 5767 13923
rect 5767 13889 5776 13923
rect 5724 13880 5776 13889
rect 5816 13923 5868 13932
rect 5816 13889 5825 13923
rect 5825 13889 5859 13923
rect 5859 13889 5868 13923
rect 5816 13880 5868 13889
rect 8300 13948 8352 14000
rect 7472 13923 7524 13932
rect 7472 13889 7481 13923
rect 7481 13889 7515 13923
rect 7515 13889 7524 13923
rect 7472 13880 7524 13889
rect 9128 13948 9180 14000
rect 9864 13948 9916 14000
rect 8484 13923 8536 13932
rect 8484 13889 8493 13923
rect 8493 13889 8527 13923
rect 8527 13889 8536 13923
rect 8484 13880 8536 13889
rect 8576 13880 8628 13932
rect 8944 13923 8996 13932
rect 8944 13889 8953 13923
rect 8953 13889 8987 13923
rect 8987 13889 8996 13923
rect 8944 13880 8996 13889
rect 9496 13923 9548 13932
rect 9496 13889 9505 13923
rect 9505 13889 9539 13923
rect 9539 13889 9548 13923
rect 9496 13880 9548 13889
rect 7564 13855 7616 13864
rect 7564 13821 7573 13855
rect 7573 13821 7607 13855
rect 7607 13821 7616 13855
rect 7564 13812 7616 13821
rect 7104 13744 7156 13796
rect 8484 13744 8536 13796
rect 9036 13744 9088 13796
rect 11060 13880 11112 13932
rect 16856 14016 16908 14068
rect 14372 13991 14424 14000
rect 14372 13957 14381 13991
rect 14381 13957 14415 13991
rect 14415 13957 14424 13991
rect 14372 13948 14424 13957
rect 12900 13880 12952 13932
rect 14096 13923 14148 13932
rect 14096 13889 14105 13923
rect 14105 13889 14139 13923
rect 14139 13889 14148 13923
rect 14096 13880 14148 13889
rect 15476 13880 15528 13932
rect 16764 13880 16816 13932
rect 11152 13812 11204 13864
rect 11244 13855 11296 13864
rect 11244 13821 11253 13855
rect 11253 13821 11287 13855
rect 11287 13821 11296 13855
rect 11244 13812 11296 13821
rect 11980 13855 12032 13864
rect 11980 13821 11989 13855
rect 11989 13821 12023 13855
rect 12023 13821 12032 13855
rect 11980 13812 12032 13821
rect 12072 13812 12124 13864
rect 12624 13812 12676 13864
rect 15108 13812 15160 13864
rect 15844 13855 15896 13864
rect 15844 13821 15853 13855
rect 15853 13821 15887 13855
rect 15887 13821 15896 13855
rect 15844 13812 15896 13821
rect 3976 13719 4028 13728
rect 3976 13685 3985 13719
rect 3985 13685 4019 13719
rect 4019 13685 4028 13719
rect 3976 13676 4028 13685
rect 6460 13676 6512 13728
rect 8760 13719 8812 13728
rect 8760 13685 8769 13719
rect 8769 13685 8803 13719
rect 8803 13685 8812 13719
rect 8760 13676 8812 13685
rect 10508 13676 10560 13728
rect 10876 13676 10928 13728
rect 15384 13744 15436 13796
rect 13360 13676 13412 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 12214 13574 12266 13626
rect 12278 13574 12330 13626
rect 12342 13574 12394 13626
rect 12406 13574 12458 13626
rect 12470 13574 12522 13626
rect 20214 13574 20266 13626
rect 20278 13574 20330 13626
rect 20342 13574 20394 13626
rect 20406 13574 20458 13626
rect 20470 13574 20522 13626
rect 2964 13515 3016 13524
rect 2964 13481 2973 13515
rect 2973 13481 3007 13515
rect 3007 13481 3016 13515
rect 2964 13472 3016 13481
rect 7472 13472 7524 13524
rect 8576 13472 8628 13524
rect 12072 13472 12124 13524
rect 14188 13472 14240 13524
rect 15752 13472 15804 13524
rect 16028 13472 16080 13524
rect 4620 13404 4672 13456
rect 3332 13336 3384 13388
rect 3240 13268 3292 13320
rect 3884 13336 3936 13388
rect 4804 13336 4856 13388
rect 3608 13268 3660 13320
rect 4712 13311 4764 13320
rect 4712 13277 4721 13311
rect 4721 13277 4755 13311
rect 4755 13277 4764 13311
rect 4712 13268 4764 13277
rect 5264 13268 5316 13320
rect 5356 13311 5408 13320
rect 5356 13277 5365 13311
rect 5365 13277 5399 13311
rect 5399 13277 5408 13311
rect 5356 13268 5408 13277
rect 5540 13311 5592 13320
rect 5540 13277 5549 13311
rect 5549 13277 5583 13311
rect 5583 13277 5592 13311
rect 5540 13268 5592 13277
rect 7288 13336 7340 13388
rect 6276 13268 6328 13320
rect 6368 13311 6420 13320
rect 6368 13277 6377 13311
rect 6377 13277 6411 13311
rect 6411 13277 6420 13311
rect 6368 13268 6420 13277
rect 6460 13311 6512 13320
rect 6460 13277 6469 13311
rect 6469 13277 6503 13311
rect 6503 13277 6512 13311
rect 6460 13268 6512 13277
rect 7104 13268 7156 13320
rect 8760 13336 8812 13388
rect 10416 13336 10468 13388
rect 12808 13336 12860 13388
rect 13268 13379 13320 13388
rect 13268 13345 13277 13379
rect 13277 13345 13311 13379
rect 13311 13345 13320 13379
rect 13268 13336 13320 13345
rect 14096 13336 14148 13388
rect 14464 13379 14516 13388
rect 14464 13345 14473 13379
rect 14473 13345 14507 13379
rect 14507 13345 14516 13379
rect 14464 13336 14516 13345
rect 6736 13200 6788 13252
rect 7012 13243 7064 13252
rect 7012 13209 7021 13243
rect 7021 13209 7055 13243
rect 7055 13209 7064 13243
rect 7012 13200 7064 13209
rect 7564 13200 7616 13252
rect 8484 13268 8536 13320
rect 9220 13311 9272 13320
rect 9220 13277 9229 13311
rect 9229 13277 9263 13311
rect 9263 13277 9272 13311
rect 9220 13268 9272 13277
rect 9588 13268 9640 13320
rect 9680 13311 9732 13320
rect 9680 13277 9689 13311
rect 9689 13277 9723 13311
rect 9723 13277 9732 13311
rect 9680 13268 9732 13277
rect 9864 13311 9916 13320
rect 9864 13277 9873 13311
rect 9873 13277 9907 13311
rect 9907 13277 9916 13311
rect 9864 13268 9916 13277
rect 13360 13311 13412 13320
rect 13360 13277 13369 13311
rect 13369 13277 13403 13311
rect 13403 13277 13412 13311
rect 13360 13268 13412 13277
rect 16764 13268 16816 13320
rect 15016 13200 15068 13252
rect 8214 13030 8266 13082
rect 8278 13030 8330 13082
rect 8342 13030 8394 13082
rect 8406 13030 8458 13082
rect 8470 13030 8522 13082
rect 16214 13030 16266 13082
rect 16278 13030 16330 13082
rect 16342 13030 16394 13082
rect 16406 13030 16458 13082
rect 16470 13030 16522 13082
rect 24214 13030 24266 13082
rect 24278 13030 24330 13082
rect 24342 13030 24394 13082
rect 24406 13030 24458 13082
rect 24470 13030 24522 13082
rect 8852 12971 8904 12980
rect 8852 12937 8861 12971
rect 8861 12937 8895 12971
rect 8895 12937 8904 12971
rect 8852 12928 8904 12937
rect 9220 12928 9272 12980
rect 10508 12971 10560 12980
rect 10508 12937 10517 12971
rect 10517 12937 10551 12971
rect 10551 12937 10560 12971
rect 10508 12928 10560 12937
rect 10784 12928 10836 12980
rect 11152 12928 11204 12980
rect 15016 12971 15068 12980
rect 15016 12937 15025 12971
rect 15025 12937 15059 12971
rect 15059 12937 15068 12971
rect 15016 12928 15068 12937
rect 15476 12971 15528 12980
rect 15476 12937 15485 12971
rect 15485 12937 15519 12971
rect 15519 12937 15528 12971
rect 15476 12928 15528 12937
rect 3608 12792 3660 12844
rect 4160 12792 4212 12844
rect 5356 12860 5408 12912
rect 4712 12792 4764 12844
rect 5264 12835 5316 12844
rect 5264 12801 5273 12835
rect 5273 12801 5307 12835
rect 5307 12801 5316 12835
rect 5264 12792 5316 12801
rect 5540 12792 5592 12844
rect 3884 12724 3936 12776
rect 4620 12724 4672 12776
rect 6276 12792 6328 12844
rect 6736 12860 6788 12912
rect 9404 12860 9456 12912
rect 10048 12860 10100 12912
rect 11060 12860 11112 12912
rect 7012 12724 7064 12776
rect 9680 12792 9732 12844
rect 9864 12792 9916 12844
rect 10876 12792 10928 12844
rect 9496 12656 9548 12708
rect 14832 12724 14884 12776
rect 15016 12792 15068 12844
rect 16028 12860 16080 12912
rect 17868 12792 17920 12844
rect 11244 12656 11296 12708
rect 8576 12588 8628 12640
rect 16672 12588 16724 12640
rect 16948 12588 17000 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 12214 12486 12266 12538
rect 12278 12486 12330 12538
rect 12342 12486 12394 12538
rect 12406 12486 12458 12538
rect 12470 12486 12522 12538
rect 20214 12486 20266 12538
rect 20278 12486 20330 12538
rect 20342 12486 20394 12538
rect 20406 12486 20458 12538
rect 20470 12486 20522 12538
rect 10876 12384 10928 12436
rect 7012 12316 7064 12368
rect 9772 12316 9824 12368
rect 10140 12316 10192 12368
rect 16764 12384 16816 12436
rect 18236 12384 18288 12436
rect 4804 12248 4856 12300
rect 11796 12248 11848 12300
rect 15568 12248 15620 12300
rect 16764 12248 16816 12300
rect 16856 12248 16908 12300
rect 17500 12291 17552 12300
rect 17500 12257 17509 12291
rect 17509 12257 17543 12291
rect 17543 12257 17552 12291
rect 17500 12248 17552 12257
rect 19616 12248 19668 12300
rect 2412 12180 2464 12232
rect 2688 12223 2740 12232
rect 2688 12189 2697 12223
rect 2697 12189 2731 12223
rect 2731 12189 2740 12223
rect 2688 12180 2740 12189
rect 3424 12180 3476 12232
rect 4896 12112 4948 12164
rect 6000 12180 6052 12232
rect 9680 12223 9732 12232
rect 9680 12189 9689 12223
rect 9689 12189 9723 12223
rect 9723 12189 9732 12223
rect 9680 12180 9732 12189
rect 6276 12112 6328 12164
rect 11244 12223 11296 12232
rect 11244 12189 11253 12223
rect 11253 12189 11287 12223
rect 11287 12189 11296 12223
rect 11244 12180 11296 12189
rect 11520 12223 11572 12232
rect 11520 12189 11529 12223
rect 11529 12189 11563 12223
rect 11563 12189 11572 12223
rect 11520 12180 11572 12189
rect 13636 12223 13688 12232
rect 13636 12189 13645 12223
rect 13645 12189 13679 12223
rect 13679 12189 13688 12223
rect 13636 12180 13688 12189
rect 14832 12223 14884 12232
rect 14832 12189 14841 12223
rect 14841 12189 14875 12223
rect 14875 12189 14884 12223
rect 14832 12180 14884 12189
rect 15016 12223 15068 12232
rect 15016 12189 15025 12223
rect 15025 12189 15059 12223
rect 15059 12189 15068 12223
rect 15016 12180 15068 12189
rect 2596 12087 2648 12096
rect 2596 12053 2605 12087
rect 2605 12053 2639 12087
rect 2639 12053 2648 12087
rect 2596 12044 2648 12053
rect 3976 12087 4028 12096
rect 3976 12053 3985 12087
rect 3985 12053 4019 12087
rect 4019 12053 4028 12087
rect 3976 12044 4028 12053
rect 5540 12044 5592 12096
rect 5816 12087 5868 12096
rect 5816 12053 5825 12087
rect 5825 12053 5859 12087
rect 5859 12053 5868 12087
rect 5816 12044 5868 12053
rect 9772 12087 9824 12096
rect 9772 12053 9781 12087
rect 9781 12053 9815 12087
rect 9815 12053 9824 12087
rect 9772 12044 9824 12053
rect 16948 12112 17000 12164
rect 17224 12155 17276 12164
rect 17224 12121 17233 12155
rect 17233 12121 17267 12155
rect 17267 12121 17276 12155
rect 17224 12112 17276 12121
rect 11704 12087 11756 12096
rect 11704 12053 11713 12087
rect 11713 12053 11747 12087
rect 11747 12053 11756 12087
rect 11704 12044 11756 12053
rect 14924 12087 14976 12096
rect 14924 12053 14933 12087
rect 14933 12053 14967 12087
rect 14967 12053 14976 12087
rect 14924 12044 14976 12053
rect 16580 12044 16632 12096
rect 16856 12044 16908 12096
rect 18236 12223 18288 12232
rect 18236 12189 18245 12223
rect 18245 12189 18279 12223
rect 18279 12189 18288 12223
rect 18236 12180 18288 12189
rect 17868 12112 17920 12164
rect 18512 12180 18564 12232
rect 19524 12112 19576 12164
rect 18328 12087 18380 12096
rect 18328 12053 18337 12087
rect 18337 12053 18371 12087
rect 18371 12053 18380 12087
rect 18328 12044 18380 12053
rect 20996 12044 21048 12096
rect 8214 11942 8266 11994
rect 8278 11942 8330 11994
rect 8342 11942 8394 11994
rect 8406 11942 8458 11994
rect 8470 11942 8522 11994
rect 16214 11942 16266 11994
rect 16278 11942 16330 11994
rect 16342 11942 16394 11994
rect 16406 11942 16458 11994
rect 16470 11942 16522 11994
rect 24214 11942 24266 11994
rect 24278 11942 24330 11994
rect 24342 11942 24394 11994
rect 24406 11942 24458 11994
rect 24470 11942 24522 11994
rect 8576 11840 8628 11892
rect 10048 11840 10100 11892
rect 10692 11883 10744 11892
rect 10692 11849 10701 11883
rect 10701 11849 10735 11883
rect 10735 11849 10744 11883
rect 10692 11840 10744 11849
rect 11244 11883 11296 11892
rect 11244 11849 11253 11883
rect 11253 11849 11287 11883
rect 11287 11849 11296 11883
rect 11244 11840 11296 11849
rect 11796 11883 11848 11892
rect 11796 11849 11805 11883
rect 11805 11849 11839 11883
rect 11839 11849 11848 11883
rect 11796 11840 11848 11849
rect 13820 11840 13872 11892
rect 14004 11840 14056 11892
rect 14280 11840 14332 11892
rect 17224 11883 17276 11892
rect 17224 11849 17233 11883
rect 17233 11849 17267 11883
rect 17267 11849 17276 11883
rect 17224 11840 17276 11849
rect 2596 11772 2648 11824
rect 5724 11772 5776 11824
rect 5816 11815 5868 11824
rect 5816 11781 5825 11815
rect 5825 11781 5859 11815
rect 5859 11781 5868 11815
rect 5816 11772 5868 11781
rect 9772 11772 9824 11824
rect 3976 11747 4028 11756
rect 3976 11713 3984 11747
rect 3984 11713 4018 11747
rect 4018 11713 4028 11747
rect 3976 11704 4028 11713
rect 4528 11704 4580 11756
rect 6920 11704 6972 11756
rect 7840 11704 7892 11756
rect 10324 11704 10376 11756
rect 14924 11772 14976 11824
rect 1492 11636 1544 11688
rect 1952 11679 2004 11688
rect 1952 11645 1961 11679
rect 1961 11645 1995 11679
rect 1995 11645 2004 11679
rect 1952 11636 2004 11645
rect 2412 11636 2464 11688
rect 6828 11636 6880 11688
rect 4620 11568 4672 11620
rect 6736 11568 6788 11620
rect 11428 11568 11480 11620
rect 3424 11543 3476 11552
rect 3424 11509 3433 11543
rect 3433 11509 3467 11543
rect 3467 11509 3476 11543
rect 3424 11500 3476 11509
rect 4068 11500 4120 11552
rect 9956 11500 10008 11552
rect 12808 11568 12860 11620
rect 13360 11568 13412 11620
rect 18328 11772 18380 11824
rect 16580 11704 16632 11756
rect 16764 11747 16816 11756
rect 16764 11713 16773 11747
rect 16773 11713 16807 11747
rect 16807 11713 16816 11747
rect 16764 11704 16816 11713
rect 17500 11704 17552 11756
rect 20996 11704 21048 11756
rect 16028 11568 16080 11620
rect 18052 11679 18104 11688
rect 18052 11645 18061 11679
rect 18061 11645 18095 11679
rect 18095 11645 18104 11679
rect 18052 11636 18104 11645
rect 19984 11636 20036 11688
rect 19064 11568 19116 11620
rect 22652 11568 22704 11620
rect 15108 11543 15160 11552
rect 15108 11509 15117 11543
rect 15117 11509 15151 11543
rect 15151 11509 15160 11543
rect 15108 11500 15160 11509
rect 16948 11543 17000 11552
rect 16948 11509 16957 11543
rect 16957 11509 16991 11543
rect 16991 11509 17000 11543
rect 16948 11500 17000 11509
rect 19800 11543 19852 11552
rect 19800 11509 19809 11543
rect 19809 11509 19843 11543
rect 19843 11509 19852 11543
rect 19800 11500 19852 11509
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 12214 11398 12266 11450
rect 12278 11398 12330 11450
rect 12342 11398 12394 11450
rect 12406 11398 12458 11450
rect 12470 11398 12522 11450
rect 20214 11398 20266 11450
rect 20278 11398 20330 11450
rect 20342 11398 20394 11450
rect 20406 11398 20458 11450
rect 20470 11398 20522 11450
rect 1952 11296 2004 11348
rect 3976 11228 4028 11280
rect 3332 11203 3384 11212
rect 3332 11169 3341 11203
rect 3341 11169 3375 11203
rect 3375 11169 3384 11203
rect 3332 11160 3384 11169
rect 3424 11092 3476 11144
rect 3976 11092 4028 11144
rect 4804 11339 4856 11348
rect 4804 11305 4813 11339
rect 4813 11305 4847 11339
rect 4847 11305 4856 11339
rect 4804 11296 4856 11305
rect 6000 11339 6052 11348
rect 6000 11305 6009 11339
rect 6009 11305 6043 11339
rect 6043 11305 6052 11339
rect 6000 11296 6052 11305
rect 6276 11339 6328 11348
rect 6276 11305 6285 11339
rect 6285 11305 6319 11339
rect 6319 11305 6328 11339
rect 6276 11296 6328 11305
rect 9956 11339 10008 11348
rect 9956 11305 9986 11339
rect 9986 11305 10008 11339
rect 9956 11296 10008 11305
rect 11428 11339 11480 11348
rect 11428 11305 11437 11339
rect 11437 11305 11471 11339
rect 11471 11305 11480 11339
rect 11428 11296 11480 11305
rect 11704 11296 11756 11348
rect 12164 11296 12216 11348
rect 14280 11296 14332 11348
rect 14832 11339 14884 11348
rect 14832 11305 14841 11339
rect 14841 11305 14875 11339
rect 14875 11305 14884 11339
rect 14832 11296 14884 11305
rect 18052 11296 18104 11348
rect 19524 11339 19576 11348
rect 19524 11305 19533 11339
rect 19533 11305 19567 11339
rect 19567 11305 19576 11339
rect 19524 11296 19576 11305
rect 22284 11296 22336 11348
rect 5540 11203 5592 11212
rect 5540 11169 5549 11203
rect 5549 11169 5583 11203
rect 5583 11169 5592 11203
rect 5540 11160 5592 11169
rect 5724 11228 5776 11280
rect 7748 11228 7800 11280
rect 7840 11228 7892 11280
rect 15568 11228 15620 11280
rect 7380 11160 7432 11212
rect 10416 11160 10468 11212
rect 14004 11160 14056 11212
rect 16948 11203 17000 11212
rect 16948 11169 16957 11203
rect 16957 11169 16991 11203
rect 16991 11169 17000 11203
rect 16948 11160 17000 11169
rect 17500 11160 17552 11212
rect 4068 11024 4120 11076
rect 6552 11135 6604 11144
rect 6552 11101 6561 11135
rect 6561 11101 6595 11135
rect 6595 11101 6604 11135
rect 6552 11092 6604 11101
rect 6828 11135 6880 11144
rect 6828 11101 6837 11135
rect 6837 11101 6871 11135
rect 6871 11101 6880 11135
rect 6828 11092 6880 11101
rect 7012 11135 7064 11144
rect 7012 11101 7021 11135
rect 7021 11101 7055 11135
rect 7055 11101 7064 11135
rect 7012 11092 7064 11101
rect 7932 11092 7984 11144
rect 9036 11092 9088 11144
rect 3240 10999 3292 11008
rect 3240 10965 3249 10999
rect 3249 10965 3283 10999
rect 3283 10965 3292 10999
rect 3240 10956 3292 10965
rect 4712 11024 4764 11076
rect 4804 10956 4856 11008
rect 8116 10999 8168 11008
rect 8116 10965 8125 10999
rect 8125 10965 8159 10999
rect 8159 10965 8168 10999
rect 8116 10956 8168 10965
rect 9312 11067 9364 11076
rect 9312 11033 9321 11067
rect 9321 11033 9355 11067
rect 9355 11033 9364 11067
rect 9312 11024 9364 11033
rect 11060 11092 11112 11144
rect 13636 11092 13688 11144
rect 19984 11160 20036 11212
rect 19064 11092 19116 11144
rect 19800 11092 19852 11144
rect 20996 11203 21048 11212
rect 20996 11169 21005 11203
rect 21005 11169 21039 11203
rect 21039 11169 21048 11203
rect 20996 11160 21048 11169
rect 9864 10956 9916 11008
rect 12624 11024 12676 11076
rect 13820 11024 13872 11076
rect 14740 11067 14792 11076
rect 14740 11033 14749 11067
rect 14749 11033 14783 11067
rect 14783 11033 14792 11067
rect 14740 11024 14792 11033
rect 16672 11024 16724 11076
rect 18052 11024 18104 11076
rect 22652 11203 22704 11212
rect 22652 11169 22661 11203
rect 22661 11169 22695 11203
rect 22695 11169 22704 11203
rect 22652 11160 22704 11169
rect 23388 11160 23440 11212
rect 10048 10956 10100 11008
rect 11244 10956 11296 11008
rect 12716 10956 12768 11008
rect 13728 10956 13780 11008
rect 15476 10999 15528 11008
rect 15476 10965 15485 10999
rect 15485 10965 15519 10999
rect 15519 10965 15528 10999
rect 15476 10956 15528 10965
rect 18236 10956 18288 11008
rect 23848 11024 23900 11076
rect 20076 10956 20128 11008
rect 21916 10956 21968 11008
rect 8214 10854 8266 10906
rect 8278 10854 8330 10906
rect 8342 10854 8394 10906
rect 8406 10854 8458 10906
rect 8470 10854 8522 10906
rect 16214 10854 16266 10906
rect 16278 10854 16330 10906
rect 16342 10854 16394 10906
rect 16406 10854 16458 10906
rect 16470 10854 16522 10906
rect 24214 10854 24266 10906
rect 24278 10854 24330 10906
rect 24342 10854 24394 10906
rect 24406 10854 24458 10906
rect 24470 10854 24522 10906
rect 3240 10752 3292 10804
rect 4712 10795 4764 10804
rect 4712 10761 4721 10795
rect 4721 10761 4755 10795
rect 4755 10761 4764 10795
rect 4712 10752 4764 10761
rect 4988 10752 5040 10804
rect 6920 10752 6972 10804
rect 7380 10795 7432 10804
rect 7380 10761 7389 10795
rect 7389 10761 7423 10795
rect 7423 10761 7432 10795
rect 7380 10752 7432 10761
rect 1308 10684 1360 10736
rect 2412 10659 2464 10668
rect 2412 10625 2421 10659
rect 2421 10625 2455 10659
rect 2455 10625 2464 10659
rect 2412 10616 2464 10625
rect 2688 10616 2740 10668
rect 6644 10684 6696 10736
rect 3976 10616 4028 10668
rect 4620 10616 4672 10668
rect 4068 10548 4120 10600
rect 3240 10480 3292 10532
rect 5540 10548 5592 10600
rect 5816 10659 5868 10668
rect 5816 10625 5825 10659
rect 5825 10625 5859 10659
rect 5859 10625 5868 10659
rect 5816 10616 5868 10625
rect 6092 10616 6144 10668
rect 8024 10752 8076 10804
rect 8116 10727 8168 10736
rect 8116 10693 8125 10727
rect 8125 10693 8159 10727
rect 8159 10693 8168 10727
rect 8116 10684 8168 10693
rect 10324 10752 10376 10804
rect 11428 10752 11480 10804
rect 11520 10752 11572 10804
rect 12716 10752 12768 10804
rect 13360 10795 13412 10804
rect 13360 10761 13369 10795
rect 13369 10761 13403 10795
rect 13403 10761 13412 10795
rect 13360 10752 13412 10761
rect 12348 10684 12400 10736
rect 12900 10684 12952 10736
rect 7840 10659 7892 10668
rect 7840 10625 7849 10659
rect 7849 10625 7883 10659
rect 7883 10625 7892 10659
rect 7840 10616 7892 10625
rect 9864 10659 9916 10668
rect 9864 10625 9873 10659
rect 9873 10625 9907 10659
rect 9907 10625 9916 10659
rect 9864 10616 9916 10625
rect 10048 10659 10100 10668
rect 10048 10625 10057 10659
rect 10057 10625 10091 10659
rect 10091 10625 10100 10659
rect 10048 10616 10100 10625
rect 10784 10659 10836 10668
rect 10784 10625 10793 10659
rect 10793 10625 10827 10659
rect 10827 10625 10836 10659
rect 10784 10616 10836 10625
rect 11336 10616 11388 10668
rect 6184 10548 6236 10600
rect 6460 10591 6512 10600
rect 6460 10557 6469 10591
rect 6469 10557 6503 10591
rect 6503 10557 6512 10591
rect 6460 10548 6512 10557
rect 10324 10548 10376 10600
rect 12716 10616 12768 10668
rect 13728 10752 13780 10804
rect 16764 10752 16816 10804
rect 15108 10684 15160 10736
rect 15292 10684 15344 10736
rect 18052 10684 18104 10736
rect 14924 10616 14976 10668
rect 15476 10616 15528 10668
rect 16120 10616 16172 10668
rect 16764 10659 16816 10668
rect 16764 10625 16773 10659
rect 16773 10625 16807 10659
rect 16807 10625 16816 10659
rect 16764 10616 16816 10625
rect 17500 10616 17552 10668
rect 19156 10616 19208 10668
rect 22560 10752 22612 10804
rect 22284 10727 22336 10736
rect 22284 10693 22293 10727
rect 22293 10693 22327 10727
rect 22327 10693 22336 10727
rect 22284 10684 22336 10693
rect 22744 10684 22796 10736
rect 21180 10659 21232 10668
rect 21180 10625 21189 10659
rect 21189 10625 21223 10659
rect 21223 10625 21232 10659
rect 21180 10616 21232 10625
rect 21732 10616 21784 10668
rect 6552 10523 6604 10532
rect 2504 10412 2556 10464
rect 6552 10489 6561 10523
rect 6561 10489 6595 10523
rect 6595 10489 6604 10523
rect 6552 10480 6604 10489
rect 9496 10480 9548 10532
rect 12164 10480 12216 10532
rect 18788 10548 18840 10600
rect 19616 10548 19668 10600
rect 4896 10412 4948 10464
rect 5448 10412 5500 10464
rect 5632 10455 5684 10464
rect 5632 10421 5641 10455
rect 5641 10421 5675 10455
rect 5675 10421 5684 10455
rect 5632 10412 5684 10421
rect 5724 10412 5776 10464
rect 6368 10412 6420 10464
rect 9404 10412 9456 10464
rect 10784 10412 10836 10464
rect 11152 10412 11204 10464
rect 12348 10412 12400 10464
rect 16028 10480 16080 10532
rect 14464 10412 14516 10464
rect 15200 10412 15252 10464
rect 16948 10455 17000 10464
rect 16948 10421 16957 10455
rect 16957 10421 16991 10455
rect 16991 10421 17000 10455
rect 16948 10412 17000 10421
rect 18696 10412 18748 10464
rect 21180 10455 21232 10464
rect 21180 10421 21189 10455
rect 21189 10421 21223 10455
rect 21223 10421 21232 10455
rect 21180 10412 21232 10421
rect 23848 10412 23900 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 12214 10310 12266 10362
rect 12278 10310 12330 10362
rect 12342 10310 12394 10362
rect 12406 10310 12458 10362
rect 12470 10310 12522 10362
rect 20214 10310 20266 10362
rect 20278 10310 20330 10362
rect 20342 10310 20394 10362
rect 20406 10310 20458 10362
rect 20470 10310 20522 10362
rect 6460 10208 6512 10260
rect 6920 10251 6972 10260
rect 6920 10217 6929 10251
rect 6929 10217 6963 10251
rect 6963 10217 6972 10251
rect 6920 10208 6972 10217
rect 7932 10251 7984 10260
rect 7932 10217 7941 10251
rect 7941 10217 7975 10251
rect 7975 10217 7984 10251
rect 7932 10208 7984 10217
rect 9036 10251 9088 10260
rect 9036 10217 9045 10251
rect 9045 10217 9079 10251
rect 9079 10217 9088 10251
rect 9036 10208 9088 10217
rect 9220 10208 9272 10260
rect 3976 10140 4028 10192
rect 4252 10072 4304 10124
rect 1492 10047 1544 10056
rect 1492 10013 1501 10047
rect 1501 10013 1535 10047
rect 1535 10013 1544 10047
rect 1492 10004 1544 10013
rect 1768 9979 1820 9988
rect 1768 9945 1777 9979
rect 1777 9945 1811 9979
rect 1811 9945 1820 9979
rect 1768 9936 1820 9945
rect 2504 9936 2556 9988
rect 4160 9936 4212 9988
rect 4436 9936 4488 9988
rect 5724 10140 5776 10192
rect 6092 10072 6144 10124
rect 6460 10072 6512 10124
rect 10324 10140 10376 10192
rect 12624 10251 12676 10260
rect 12624 10217 12633 10251
rect 12633 10217 12667 10251
rect 12667 10217 12676 10251
rect 12624 10208 12676 10217
rect 14924 10251 14976 10260
rect 14924 10217 14933 10251
rect 14933 10217 14967 10251
rect 14967 10217 14976 10251
rect 14924 10208 14976 10217
rect 16764 10208 16816 10260
rect 19156 10208 19208 10260
rect 22744 10251 22796 10260
rect 22744 10217 22753 10251
rect 22753 10217 22787 10251
rect 22787 10217 22796 10251
rect 22744 10208 22796 10217
rect 15292 10140 15344 10192
rect 5448 10004 5500 10056
rect 5816 10004 5868 10056
rect 5908 10047 5960 10056
rect 5908 10013 5917 10047
rect 5917 10013 5951 10047
rect 5951 10013 5960 10047
rect 5908 10004 5960 10013
rect 6184 10047 6236 10056
rect 6184 10013 6193 10047
rect 6193 10013 6227 10047
rect 6227 10013 6236 10047
rect 6184 10004 6236 10013
rect 6276 10047 6328 10056
rect 6276 10013 6286 10047
rect 6286 10013 6320 10047
rect 6320 10013 6328 10047
rect 6276 10004 6328 10013
rect 6920 10004 6972 10056
rect 9496 10115 9548 10124
rect 9496 10081 9505 10115
rect 9505 10081 9539 10115
rect 9539 10081 9548 10115
rect 9496 10072 9548 10081
rect 9680 10115 9732 10124
rect 9680 10081 9689 10115
rect 9689 10081 9723 10115
rect 9723 10081 9732 10115
rect 9680 10072 9732 10081
rect 10416 10115 10468 10124
rect 10416 10081 10425 10115
rect 10425 10081 10459 10115
rect 10459 10081 10468 10115
rect 10416 10072 10468 10081
rect 11244 10072 11296 10124
rect 7564 10004 7616 10056
rect 7932 10004 7984 10056
rect 12900 10072 12952 10124
rect 15108 10072 15160 10124
rect 16580 10072 16632 10124
rect 18236 10115 18288 10124
rect 18236 10081 18245 10115
rect 18245 10081 18279 10115
rect 18279 10081 18288 10115
rect 18236 10072 18288 10081
rect 5540 9936 5592 9988
rect 6092 9936 6144 9988
rect 3240 9911 3292 9920
rect 3240 9877 3249 9911
rect 3249 9877 3283 9911
rect 3283 9877 3292 9911
rect 3240 9868 3292 9877
rect 5356 9868 5408 9920
rect 6552 9868 6604 9920
rect 6644 9868 6696 9920
rect 8760 9936 8812 9988
rect 10692 9979 10744 9988
rect 10692 9945 10701 9979
rect 10701 9945 10735 9979
rect 10735 9945 10744 9979
rect 10692 9936 10744 9945
rect 11980 9936 12032 9988
rect 12716 10004 12768 10056
rect 9220 9868 9272 9920
rect 11704 9868 11756 9920
rect 12164 9911 12216 9920
rect 12164 9877 12173 9911
rect 12173 9877 12207 9911
rect 12207 9877 12216 9911
rect 12164 9868 12216 9877
rect 13084 9868 13136 9920
rect 15384 9936 15436 9988
rect 15292 9911 15344 9920
rect 15292 9877 15301 9911
rect 15301 9877 15335 9911
rect 15335 9877 15344 9911
rect 15292 9868 15344 9877
rect 16028 10047 16080 10056
rect 16028 10013 16037 10047
rect 16037 10013 16071 10047
rect 16071 10013 16080 10047
rect 16028 10004 16080 10013
rect 16120 10004 16172 10056
rect 18696 10004 18748 10056
rect 19156 10004 19208 10056
rect 19616 10072 19668 10124
rect 23388 10140 23440 10192
rect 21088 10072 21140 10124
rect 21456 10072 21508 10124
rect 19524 10047 19576 10056
rect 19524 10013 19533 10047
rect 19533 10013 19567 10047
rect 19567 10013 19576 10047
rect 19524 10004 19576 10013
rect 22560 10047 22612 10056
rect 22560 10013 22569 10047
rect 22569 10013 22603 10047
rect 22603 10013 22612 10047
rect 22560 10004 22612 10013
rect 17776 9936 17828 9988
rect 18972 9868 19024 9920
rect 20076 9936 20128 9988
rect 21180 9936 21232 9988
rect 24124 10004 24176 10056
rect 24768 9936 24820 9988
rect 21916 9911 21968 9920
rect 21916 9877 21925 9911
rect 21925 9877 21959 9911
rect 21959 9877 21968 9911
rect 21916 9868 21968 9877
rect 22744 9868 22796 9920
rect 8214 9766 8266 9818
rect 8278 9766 8330 9818
rect 8342 9766 8394 9818
rect 8406 9766 8458 9818
rect 8470 9766 8522 9818
rect 16214 9766 16266 9818
rect 16278 9766 16330 9818
rect 16342 9766 16394 9818
rect 16406 9766 16458 9818
rect 16470 9766 16522 9818
rect 24214 9766 24266 9818
rect 24278 9766 24330 9818
rect 24342 9766 24394 9818
rect 24406 9766 24458 9818
rect 24470 9766 24522 9818
rect 1768 9664 1820 9716
rect 3240 9664 3292 9716
rect 5908 9664 5960 9716
rect 4252 9596 4304 9648
rect 4436 9596 4488 9648
rect 4528 9528 4580 9580
rect 3424 9460 3476 9512
rect 3976 9392 4028 9444
rect 4712 9392 4764 9444
rect 4988 9392 5040 9444
rect 4068 9324 4120 9376
rect 5356 9571 5408 9580
rect 5356 9537 5365 9571
rect 5365 9537 5399 9571
rect 5399 9537 5408 9571
rect 5356 9528 5408 9537
rect 5632 9528 5684 9580
rect 5724 9571 5776 9580
rect 5724 9537 5733 9571
rect 5733 9537 5767 9571
rect 5767 9537 5776 9571
rect 5724 9528 5776 9537
rect 6092 9639 6144 9648
rect 6092 9605 6101 9639
rect 6101 9605 6135 9639
rect 6135 9605 6144 9639
rect 6092 9596 6144 9605
rect 6552 9639 6604 9648
rect 6552 9605 6561 9639
rect 6561 9605 6595 9639
rect 6595 9605 6604 9639
rect 6552 9596 6604 9605
rect 9220 9707 9272 9716
rect 9220 9673 9229 9707
rect 9229 9673 9263 9707
rect 9263 9673 9272 9707
rect 9220 9664 9272 9673
rect 10692 9664 10744 9716
rect 15292 9664 15344 9716
rect 18788 9707 18840 9716
rect 18788 9673 18797 9707
rect 18797 9673 18831 9707
rect 18831 9673 18840 9707
rect 18788 9664 18840 9673
rect 19524 9664 19576 9716
rect 5908 9528 5960 9580
rect 6276 9528 6328 9580
rect 6736 9571 6788 9580
rect 6736 9537 6745 9571
rect 6745 9537 6779 9571
rect 6779 9537 6788 9571
rect 6736 9528 6788 9537
rect 7196 9528 7248 9580
rect 7840 9596 7892 9648
rect 9312 9596 9364 9648
rect 9864 9596 9916 9648
rect 10784 9596 10836 9648
rect 10416 9528 10468 9580
rect 10692 9571 10744 9580
rect 10692 9537 10701 9571
rect 10701 9537 10735 9571
rect 10735 9537 10744 9571
rect 10692 9528 10744 9537
rect 11704 9596 11756 9648
rect 11244 9571 11296 9580
rect 11244 9537 11253 9571
rect 11253 9537 11287 9571
rect 11287 9537 11296 9571
rect 11244 9528 11296 9537
rect 11980 9639 12032 9648
rect 11980 9605 11989 9639
rect 11989 9605 12023 9639
rect 12023 9605 12032 9639
rect 11980 9596 12032 9605
rect 14464 9639 14516 9648
rect 14464 9605 14473 9639
rect 14473 9605 14507 9639
rect 14507 9605 14516 9639
rect 14464 9596 14516 9605
rect 15476 9596 15528 9648
rect 16948 9596 17000 9648
rect 17684 9596 17736 9648
rect 22560 9664 22612 9716
rect 23480 9664 23532 9716
rect 12072 9571 12124 9580
rect 12072 9537 12081 9571
rect 12081 9537 12115 9571
rect 12115 9537 12124 9571
rect 12072 9528 12124 9537
rect 18972 9571 19024 9580
rect 18972 9537 18981 9571
rect 18981 9537 19015 9571
rect 19015 9537 19024 9571
rect 18972 9528 19024 9537
rect 19524 9571 19576 9580
rect 19524 9537 19533 9571
rect 19533 9537 19567 9571
rect 19567 9537 19576 9571
rect 19524 9528 19576 9537
rect 20904 9528 20956 9580
rect 22100 9571 22152 9580
rect 22100 9537 22109 9571
rect 22109 9537 22143 9571
rect 22143 9537 22152 9571
rect 22100 9528 22152 9537
rect 22744 9528 22796 9580
rect 23020 9571 23072 9580
rect 23020 9537 23029 9571
rect 23029 9537 23063 9571
rect 23063 9537 23072 9571
rect 23020 9528 23072 9537
rect 24400 9528 24452 9580
rect 6828 9460 6880 9512
rect 7748 9503 7800 9512
rect 7748 9469 7757 9503
rect 7757 9469 7791 9503
rect 7791 9469 7800 9503
rect 7748 9460 7800 9469
rect 13176 9460 13228 9512
rect 16672 9460 16724 9512
rect 17776 9460 17828 9512
rect 19800 9503 19852 9512
rect 19800 9469 19809 9503
rect 19809 9469 19843 9503
rect 19843 9469 19852 9503
rect 19800 9460 19852 9469
rect 21456 9460 21508 9512
rect 11060 9435 11112 9444
rect 11060 9401 11069 9435
rect 11069 9401 11103 9435
rect 11103 9401 11112 9435
rect 11060 9392 11112 9401
rect 24768 9503 24820 9512
rect 24768 9469 24777 9503
rect 24777 9469 24811 9503
rect 24811 9469 24820 9503
rect 24768 9460 24820 9469
rect 7564 9324 7616 9376
rect 9588 9324 9640 9376
rect 11520 9324 11572 9376
rect 12164 9324 12216 9376
rect 18420 9324 18472 9376
rect 22836 9324 22888 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 12214 9222 12266 9274
rect 12278 9222 12330 9274
rect 12342 9222 12394 9274
rect 12406 9222 12458 9274
rect 12470 9222 12522 9274
rect 20214 9222 20266 9274
rect 20278 9222 20330 9274
rect 20342 9222 20394 9274
rect 20406 9222 20458 9274
rect 20470 9222 20522 9274
rect 6552 9163 6604 9172
rect 6552 9129 6561 9163
rect 6561 9129 6595 9163
rect 6595 9129 6604 9163
rect 6552 9120 6604 9129
rect 6736 9120 6788 9172
rect 3976 9052 4028 9104
rect 3240 8984 3292 9036
rect 4620 9027 4672 9036
rect 4620 8993 4629 9027
rect 4629 8993 4663 9027
rect 4663 8993 4672 9027
rect 4620 8984 4672 8993
rect 2228 8959 2280 8968
rect 2228 8925 2237 8959
rect 2237 8925 2271 8959
rect 2271 8925 2280 8959
rect 2228 8916 2280 8925
rect 3608 8916 3660 8968
rect 4712 8916 4764 8968
rect 4988 8916 5040 8968
rect 11152 9120 11204 9172
rect 15476 9163 15528 9172
rect 15476 9129 15485 9163
rect 15485 9129 15519 9163
rect 15519 9129 15528 9163
rect 15476 9120 15528 9129
rect 17684 9163 17736 9172
rect 17684 9129 17693 9163
rect 17693 9129 17727 9163
rect 17727 9129 17736 9163
rect 17684 9120 17736 9129
rect 22100 9120 22152 9172
rect 24400 9120 24452 9172
rect 7840 8984 7892 9036
rect 9588 9027 9640 9036
rect 9588 8993 9597 9027
rect 9597 8993 9631 9027
rect 9631 8993 9640 9027
rect 9588 8984 9640 8993
rect 13176 8984 13228 9036
rect 14556 9027 14608 9036
rect 14556 8993 14565 9027
rect 14565 8993 14599 9027
rect 14599 8993 14608 9027
rect 14556 8984 14608 8993
rect 7104 8916 7156 8968
rect 8024 8916 8076 8968
rect 15292 8916 15344 8968
rect 15384 8916 15436 8968
rect 1768 8780 1820 8832
rect 4528 8823 4580 8832
rect 4528 8789 4537 8823
rect 4537 8789 4571 8823
rect 4571 8789 4580 8823
rect 4528 8780 4580 8789
rect 4712 8780 4764 8832
rect 4896 8780 4948 8832
rect 6000 8780 6052 8832
rect 7288 8780 7340 8832
rect 10600 8848 10652 8900
rect 11888 8848 11940 8900
rect 15660 8959 15712 8968
rect 15660 8925 15669 8959
rect 15669 8925 15703 8959
rect 15703 8925 15712 8959
rect 15660 8916 15712 8925
rect 11704 8823 11756 8832
rect 11704 8789 11713 8823
rect 11713 8789 11747 8823
rect 11747 8789 11756 8823
rect 11704 8780 11756 8789
rect 12440 8780 12492 8832
rect 16028 8848 16080 8900
rect 17224 9052 17276 9104
rect 18420 8984 18472 9036
rect 19984 9027 20036 9036
rect 19984 8993 19993 9027
rect 19993 8993 20027 9027
rect 20027 8993 20036 9027
rect 19984 8984 20036 8993
rect 22836 9027 22888 9036
rect 22836 8993 22845 9027
rect 22845 8993 22879 9027
rect 22879 8993 22888 9027
rect 22836 8984 22888 8993
rect 23112 9027 23164 9036
rect 23112 8993 23121 9027
rect 23121 8993 23155 9027
rect 23155 8993 23164 9027
rect 23112 8984 23164 8993
rect 23388 8984 23440 9036
rect 16488 8916 16540 8968
rect 14832 8823 14884 8832
rect 14832 8789 14841 8823
rect 14841 8789 14875 8823
rect 14875 8789 14884 8823
rect 14832 8780 14884 8789
rect 15476 8780 15528 8832
rect 17500 8848 17552 8900
rect 17960 8916 18012 8968
rect 21456 8916 21508 8968
rect 24124 8916 24176 8968
rect 19156 8848 19208 8900
rect 20076 8848 20128 8900
rect 21824 8848 21876 8900
rect 23480 8848 23532 8900
rect 16488 8780 16540 8832
rect 19524 8780 19576 8832
rect 20628 8823 20680 8832
rect 20628 8789 20637 8823
rect 20637 8789 20671 8823
rect 20671 8789 20680 8823
rect 20628 8780 20680 8789
rect 24124 8780 24176 8832
rect 8214 8678 8266 8730
rect 8278 8678 8330 8730
rect 8342 8678 8394 8730
rect 8406 8678 8458 8730
rect 8470 8678 8522 8730
rect 16214 8678 16266 8730
rect 16278 8678 16330 8730
rect 16342 8678 16394 8730
rect 16406 8678 16458 8730
rect 16470 8678 16522 8730
rect 24214 8678 24266 8730
rect 24278 8678 24330 8730
rect 24342 8678 24394 8730
rect 24406 8678 24458 8730
rect 24470 8678 24522 8730
rect 1308 8576 1360 8628
rect 1768 8551 1820 8560
rect 1768 8517 1777 8551
rect 1777 8517 1811 8551
rect 1811 8517 1820 8551
rect 1768 8508 1820 8517
rect 2780 8508 2832 8560
rect 3608 8619 3660 8628
rect 3608 8585 3617 8619
rect 3617 8585 3651 8619
rect 3651 8585 3660 8619
rect 3608 8576 3660 8585
rect 3884 8576 3936 8628
rect 7104 8576 7156 8628
rect 8300 8576 8352 8628
rect 10416 8619 10468 8628
rect 10416 8585 10425 8619
rect 10425 8585 10459 8619
rect 10459 8585 10468 8619
rect 10416 8576 10468 8585
rect 10600 8576 10652 8628
rect 11888 8619 11940 8628
rect 11888 8585 11897 8619
rect 11897 8585 11931 8619
rect 11931 8585 11940 8619
rect 11888 8576 11940 8585
rect 12440 8619 12492 8628
rect 12440 8585 12449 8619
rect 12449 8585 12483 8619
rect 12483 8585 12492 8619
rect 12440 8576 12492 8585
rect 5080 8508 5132 8560
rect 7380 8508 7432 8560
rect 11520 8508 11572 8560
rect 4068 8440 4120 8492
rect 1492 8415 1544 8424
rect 1492 8381 1501 8415
rect 1501 8381 1535 8415
rect 1535 8381 1544 8415
rect 1492 8372 1544 8381
rect 3240 8415 3292 8424
rect 3240 8381 3249 8415
rect 3249 8381 3283 8415
rect 3283 8381 3292 8415
rect 3240 8372 3292 8381
rect 4804 8440 4856 8492
rect 5172 8483 5224 8492
rect 5172 8449 5181 8483
rect 5181 8449 5215 8483
rect 5215 8449 5224 8483
rect 5172 8440 5224 8449
rect 4712 8415 4764 8424
rect 4712 8381 4721 8415
rect 4721 8381 4755 8415
rect 4755 8381 4764 8415
rect 4712 8372 4764 8381
rect 4896 8372 4948 8424
rect 7104 8440 7156 8492
rect 7196 8483 7248 8492
rect 7196 8449 7205 8483
rect 7205 8449 7239 8483
rect 7239 8449 7248 8483
rect 7196 8440 7248 8449
rect 6000 8415 6052 8424
rect 6000 8381 6009 8415
rect 6009 8381 6043 8415
rect 6043 8381 6052 8415
rect 6000 8372 6052 8381
rect 9680 8440 9732 8492
rect 10784 8440 10836 8492
rect 9312 8372 9364 8424
rect 9772 8415 9824 8424
rect 9772 8381 9781 8415
rect 9781 8381 9815 8415
rect 9815 8381 9824 8415
rect 9772 8372 9824 8381
rect 10600 8372 10652 8424
rect 11244 8440 11296 8492
rect 11888 8440 11940 8492
rect 11980 8483 12032 8492
rect 11980 8449 11989 8483
rect 11989 8449 12023 8483
rect 12023 8449 12032 8483
rect 11980 8440 12032 8449
rect 17224 8576 17276 8628
rect 15016 8508 15068 8560
rect 15476 8551 15528 8560
rect 15476 8517 15485 8551
rect 15485 8517 15519 8551
rect 15519 8517 15528 8551
rect 15476 8508 15528 8517
rect 17776 8619 17828 8628
rect 17776 8585 17785 8619
rect 17785 8585 17819 8619
rect 17819 8585 17828 8619
rect 17776 8576 17828 8585
rect 18696 8619 18748 8628
rect 18696 8585 18705 8619
rect 18705 8585 18739 8619
rect 18739 8585 18748 8619
rect 18696 8576 18748 8585
rect 19800 8576 19852 8628
rect 20904 8576 20956 8628
rect 21824 8576 21876 8628
rect 18972 8508 19024 8560
rect 19248 8508 19300 8560
rect 11704 8372 11756 8424
rect 17592 8440 17644 8492
rect 18788 8483 18840 8492
rect 18788 8449 18797 8483
rect 18797 8449 18831 8483
rect 18831 8449 18840 8483
rect 18788 8440 18840 8449
rect 19524 8483 19576 8492
rect 19524 8449 19533 8483
rect 19533 8449 19567 8483
rect 19567 8449 19576 8483
rect 19524 8440 19576 8449
rect 20628 8508 20680 8560
rect 4528 8304 4580 8356
rect 5540 8347 5592 8356
rect 5540 8313 5549 8347
rect 5549 8313 5583 8347
rect 5583 8313 5592 8347
rect 5540 8304 5592 8313
rect 8760 8304 8812 8356
rect 14832 8372 14884 8424
rect 16672 8372 16724 8424
rect 17500 8372 17552 8424
rect 13820 8304 13872 8356
rect 14464 8304 14516 8356
rect 19432 8304 19484 8356
rect 19616 8372 19668 8424
rect 20812 8483 20864 8492
rect 20812 8449 20821 8483
rect 20821 8449 20855 8483
rect 20855 8449 20864 8483
rect 20812 8440 20864 8449
rect 23572 8508 23624 8560
rect 21824 8440 21876 8492
rect 22008 8372 22060 8424
rect 16948 8236 17000 8288
rect 20076 8304 20128 8356
rect 23112 8440 23164 8492
rect 23664 8415 23716 8424
rect 23664 8381 23673 8415
rect 23673 8381 23707 8415
rect 23707 8381 23716 8415
rect 23664 8372 23716 8381
rect 20720 8236 20772 8288
rect 20996 8279 21048 8288
rect 20996 8245 21005 8279
rect 21005 8245 21039 8279
rect 21039 8245 21048 8279
rect 20996 8236 21048 8245
rect 22928 8236 22980 8288
rect 23480 8236 23532 8288
rect 25136 8279 25188 8288
rect 25136 8245 25145 8279
rect 25145 8245 25179 8279
rect 25179 8245 25188 8279
rect 25136 8236 25188 8245
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 12214 8134 12266 8186
rect 12278 8134 12330 8186
rect 12342 8134 12394 8186
rect 12406 8134 12458 8186
rect 12470 8134 12522 8186
rect 20214 8134 20266 8186
rect 20278 8134 20330 8186
rect 20342 8134 20394 8186
rect 20406 8134 20458 8186
rect 20470 8134 20522 8186
rect 2228 8032 2280 8084
rect 3608 8032 3660 8084
rect 4620 8032 4672 8084
rect 2780 7964 2832 8016
rect 2504 7896 2556 7948
rect 5172 7964 5224 8016
rect 6368 8032 6420 8084
rect 10692 8075 10744 8084
rect 10692 8041 10701 8075
rect 10701 8041 10735 8075
rect 10735 8041 10744 8075
rect 10692 8032 10744 8041
rect 11888 8032 11940 8084
rect 12256 8032 12308 8084
rect 14556 8032 14608 8084
rect 15016 8032 15068 8084
rect 9680 8007 9732 8016
rect 3424 7896 3476 7948
rect 9680 7973 9689 8007
rect 9689 7973 9723 8007
rect 9723 7973 9732 8007
rect 9680 7964 9732 7973
rect 2688 7828 2740 7880
rect 3240 7828 3292 7880
rect 4068 7828 4120 7880
rect 4896 7828 4948 7880
rect 4436 7692 4488 7744
rect 4896 7735 4948 7744
rect 4896 7701 4905 7735
rect 4905 7701 4939 7735
rect 4939 7701 4948 7735
rect 4896 7692 4948 7701
rect 5816 7871 5868 7880
rect 5816 7837 5825 7871
rect 5825 7837 5859 7871
rect 5859 7837 5868 7871
rect 5816 7828 5868 7837
rect 6368 7871 6420 7880
rect 6368 7837 6377 7871
rect 6377 7837 6411 7871
rect 6411 7837 6420 7871
rect 6368 7828 6420 7837
rect 8576 7896 8628 7948
rect 9772 7896 9824 7948
rect 11152 7896 11204 7948
rect 8116 7828 8168 7880
rect 8300 7871 8352 7880
rect 8300 7837 8309 7871
rect 8309 7837 8343 7871
rect 8343 7837 8352 7871
rect 8300 7828 8352 7837
rect 8668 7828 8720 7880
rect 12072 7828 12124 7880
rect 5540 7803 5592 7812
rect 5540 7769 5549 7803
rect 5549 7769 5583 7803
rect 5583 7769 5592 7803
rect 5540 7760 5592 7769
rect 6000 7760 6052 7812
rect 10140 7760 10192 7812
rect 11796 7760 11848 7812
rect 14188 7871 14240 7880
rect 14188 7837 14197 7871
rect 14197 7837 14231 7871
rect 14231 7837 14240 7871
rect 14188 7828 14240 7837
rect 14740 7828 14792 7880
rect 15200 7760 15252 7812
rect 15660 7828 15712 7880
rect 16028 7871 16080 7880
rect 16028 7837 16037 7871
rect 16037 7837 16071 7871
rect 16071 7837 16080 7871
rect 16028 7828 16080 7837
rect 18236 8032 18288 8084
rect 16948 7939 17000 7948
rect 16948 7905 16957 7939
rect 16957 7905 16991 7939
rect 16991 7905 17000 7939
rect 16948 7896 17000 7905
rect 16672 7871 16724 7880
rect 16672 7837 16681 7871
rect 16681 7837 16715 7871
rect 16715 7837 16724 7871
rect 16672 7828 16724 7837
rect 23572 8032 23624 8084
rect 23664 8032 23716 8084
rect 24032 8032 24084 8084
rect 23112 7964 23164 8016
rect 20996 7896 21048 7948
rect 22376 7896 22428 7948
rect 18972 7828 19024 7880
rect 19432 7828 19484 7880
rect 20352 7828 20404 7880
rect 23112 7871 23164 7880
rect 23112 7837 23121 7871
rect 23121 7837 23155 7871
rect 23155 7837 23164 7871
rect 23112 7828 23164 7837
rect 5724 7735 5776 7744
rect 5724 7701 5733 7735
rect 5733 7701 5767 7735
rect 5767 7701 5776 7735
rect 5724 7692 5776 7701
rect 7748 7692 7800 7744
rect 8024 7692 8076 7744
rect 8944 7692 8996 7744
rect 12900 7735 12952 7744
rect 12900 7701 12909 7735
rect 12909 7701 12943 7735
rect 12943 7701 12952 7735
rect 12900 7692 12952 7701
rect 13636 7692 13688 7744
rect 22560 7760 22612 7812
rect 23480 7828 23532 7880
rect 24768 7896 24820 7948
rect 25136 7828 25188 7880
rect 15844 7692 15896 7744
rect 17592 7692 17644 7744
rect 18880 7692 18932 7744
rect 21088 7692 21140 7744
rect 22652 7692 22704 7744
rect 8214 7590 8266 7642
rect 8278 7590 8330 7642
rect 8342 7590 8394 7642
rect 8406 7590 8458 7642
rect 8470 7590 8522 7642
rect 16214 7590 16266 7642
rect 16278 7590 16330 7642
rect 16342 7590 16394 7642
rect 16406 7590 16458 7642
rect 16470 7590 16522 7642
rect 24214 7590 24266 7642
rect 24278 7590 24330 7642
rect 24342 7590 24394 7642
rect 24406 7590 24458 7642
rect 24470 7590 24522 7642
rect 4436 7531 4488 7540
rect 4436 7497 4445 7531
rect 4445 7497 4479 7531
rect 4479 7497 4488 7531
rect 4436 7488 4488 7497
rect 5724 7488 5776 7540
rect 5816 7488 5868 7540
rect 6092 7488 6144 7540
rect 7104 7531 7156 7540
rect 7104 7497 7113 7531
rect 7113 7497 7147 7531
rect 7147 7497 7156 7531
rect 7104 7488 7156 7497
rect 1860 7352 1912 7404
rect 2504 7395 2556 7404
rect 2504 7361 2513 7395
rect 2513 7361 2547 7395
rect 2547 7361 2556 7395
rect 2504 7352 2556 7361
rect 2688 7395 2740 7404
rect 2688 7361 2697 7395
rect 2697 7361 2731 7395
rect 2731 7361 2740 7395
rect 2688 7352 2740 7361
rect 4068 7395 4120 7404
rect 4068 7361 4076 7395
rect 4076 7361 4110 7395
rect 4110 7361 4120 7395
rect 4068 7352 4120 7361
rect 4896 7420 4948 7472
rect 6276 7420 6328 7472
rect 11060 7488 11112 7540
rect 5172 7352 5224 7404
rect 8024 7463 8076 7472
rect 8024 7429 8033 7463
rect 8033 7429 8067 7463
rect 8067 7429 8076 7463
rect 8024 7420 8076 7429
rect 9588 7420 9640 7472
rect 5540 7216 5592 7268
rect 6644 7395 6696 7404
rect 6644 7361 6653 7395
rect 6653 7361 6687 7395
rect 6687 7361 6696 7395
rect 6644 7352 6696 7361
rect 7012 7395 7064 7404
rect 7012 7361 7021 7395
rect 7021 7361 7055 7395
rect 7055 7361 7064 7395
rect 7012 7352 7064 7361
rect 10140 7352 10192 7404
rect 11796 7395 11848 7404
rect 11796 7361 11805 7395
rect 11805 7361 11839 7395
rect 11839 7361 11848 7395
rect 11796 7352 11848 7361
rect 11980 7352 12032 7404
rect 13636 7488 13688 7540
rect 14188 7488 14240 7540
rect 12900 7420 12952 7472
rect 16672 7488 16724 7540
rect 15108 7420 15160 7472
rect 18880 7463 18932 7472
rect 18880 7429 18889 7463
rect 18889 7429 18923 7463
rect 18923 7429 18932 7463
rect 18880 7420 18932 7429
rect 12256 7395 12308 7404
rect 12256 7361 12265 7395
rect 12265 7361 12299 7395
rect 12299 7361 12308 7395
rect 12256 7352 12308 7361
rect 15660 7352 15712 7404
rect 16948 7395 17000 7404
rect 16948 7361 16957 7395
rect 16957 7361 16991 7395
rect 16991 7361 17000 7395
rect 16948 7352 17000 7361
rect 17776 7352 17828 7404
rect 20352 7531 20404 7540
rect 20352 7497 20361 7531
rect 20361 7497 20395 7531
rect 20395 7497 20404 7531
rect 20352 7488 20404 7497
rect 20812 7488 20864 7540
rect 21088 7531 21140 7540
rect 21088 7497 21097 7531
rect 21097 7497 21131 7531
rect 21131 7497 21140 7531
rect 21088 7488 21140 7497
rect 21916 7488 21968 7540
rect 24124 7531 24176 7540
rect 24124 7497 24133 7531
rect 24133 7497 24167 7531
rect 24167 7497 24176 7531
rect 24124 7488 24176 7497
rect 19432 7420 19484 7472
rect 19248 7352 19300 7404
rect 20076 7352 20128 7404
rect 22560 7420 22612 7472
rect 22652 7463 22704 7472
rect 22652 7429 22661 7463
rect 22661 7429 22695 7463
rect 22695 7429 22704 7463
rect 22652 7420 22704 7429
rect 22928 7420 22980 7472
rect 21824 7352 21876 7404
rect 22008 7352 22060 7404
rect 22376 7395 22428 7404
rect 22376 7361 22385 7395
rect 22385 7361 22419 7395
rect 22419 7361 22428 7395
rect 22376 7352 22428 7361
rect 24584 7395 24636 7404
rect 24584 7361 24593 7395
rect 24593 7361 24627 7395
rect 24627 7361 24636 7395
rect 24584 7352 24636 7361
rect 7196 7284 7248 7336
rect 9036 7284 9088 7336
rect 13176 7327 13228 7336
rect 13176 7293 13185 7327
rect 13185 7293 13219 7327
rect 13219 7293 13228 7327
rect 13176 7284 13228 7293
rect 13452 7327 13504 7336
rect 13452 7293 13461 7327
rect 13461 7293 13495 7327
rect 13495 7293 13504 7327
rect 13452 7284 13504 7293
rect 15384 7284 15436 7336
rect 18788 7284 18840 7336
rect 20720 7284 20772 7336
rect 24032 7284 24084 7336
rect 23940 7216 23992 7268
rect 2780 7148 2832 7200
rect 7472 7191 7524 7200
rect 7472 7157 7481 7191
rect 7481 7157 7515 7191
rect 7515 7157 7524 7191
rect 7472 7148 7524 7157
rect 9496 7191 9548 7200
rect 9496 7157 9505 7191
rect 9505 7157 9539 7191
rect 9539 7157 9548 7191
rect 9496 7148 9548 7157
rect 9956 7191 10008 7200
rect 9956 7157 9965 7191
rect 9965 7157 9999 7191
rect 9999 7157 10008 7191
rect 9956 7148 10008 7157
rect 11612 7191 11664 7200
rect 11612 7157 11621 7191
rect 11621 7157 11655 7191
rect 11655 7157 11664 7191
rect 11612 7148 11664 7157
rect 11980 7148 12032 7200
rect 14924 7191 14976 7200
rect 14924 7157 14933 7191
rect 14933 7157 14967 7191
rect 14967 7157 14976 7191
rect 14924 7148 14976 7157
rect 21916 7191 21968 7200
rect 21916 7157 21925 7191
rect 21925 7157 21959 7191
rect 21959 7157 21968 7191
rect 21916 7148 21968 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 12214 7046 12266 7098
rect 12278 7046 12330 7098
rect 12342 7046 12394 7098
rect 12406 7046 12458 7098
rect 12470 7046 12522 7098
rect 20214 7046 20266 7098
rect 20278 7046 20330 7098
rect 20342 7046 20394 7098
rect 20406 7046 20458 7098
rect 20470 7046 20522 7098
rect 4068 6944 4120 6996
rect 6000 6987 6052 6996
rect 6000 6953 6009 6987
rect 6009 6953 6043 6987
rect 6043 6953 6052 6987
rect 6000 6944 6052 6953
rect 7104 6944 7156 6996
rect 1492 6851 1544 6860
rect 1492 6817 1501 6851
rect 1501 6817 1535 6851
rect 1535 6817 1544 6851
rect 1492 6808 1544 6817
rect 5172 6808 5224 6860
rect 6644 6876 6696 6928
rect 8760 6876 8812 6928
rect 9772 6944 9824 6996
rect 11612 6944 11664 6996
rect 13452 6944 13504 6996
rect 18604 6944 18656 6996
rect 19248 6944 19300 6996
rect 19524 6944 19576 6996
rect 22376 6944 22428 6996
rect 23112 6944 23164 6996
rect 24584 6944 24636 6996
rect 9404 6876 9456 6928
rect 5540 6808 5592 6860
rect 7380 6851 7432 6860
rect 7380 6817 7389 6851
rect 7389 6817 7423 6851
rect 7423 6817 7432 6851
rect 7380 6808 7432 6817
rect 7472 6808 7524 6860
rect 1768 6715 1820 6724
rect 1768 6681 1777 6715
rect 1777 6681 1811 6715
rect 1811 6681 1820 6715
rect 1768 6672 1820 6681
rect 2780 6672 2832 6724
rect 4804 6672 4856 6724
rect 3148 6604 3200 6656
rect 4896 6604 4948 6656
rect 5632 6740 5684 6792
rect 6092 6783 6144 6792
rect 6092 6749 6101 6783
rect 6101 6749 6135 6783
rect 6135 6749 6144 6783
rect 6092 6740 6144 6749
rect 5724 6672 5776 6724
rect 7748 6783 7800 6792
rect 7748 6749 7757 6783
rect 7757 6749 7791 6783
rect 7791 6749 7800 6783
rect 7748 6740 7800 6749
rect 8668 6808 8720 6860
rect 8024 6783 8076 6792
rect 8024 6749 8033 6783
rect 8033 6749 8067 6783
rect 8067 6749 8076 6783
rect 8024 6740 8076 6749
rect 5448 6604 5500 6656
rect 6092 6604 6144 6656
rect 7104 6604 7156 6656
rect 8576 6740 8628 6792
rect 8668 6715 8720 6724
rect 8668 6681 8677 6715
rect 8677 6681 8711 6715
rect 8711 6681 8720 6715
rect 8668 6672 8720 6681
rect 9496 6808 9548 6860
rect 9588 6808 9640 6860
rect 10968 6851 11020 6860
rect 10968 6817 10977 6851
rect 10977 6817 11011 6851
rect 11011 6817 11020 6851
rect 13176 6876 13228 6928
rect 17960 6876 18012 6928
rect 18972 6876 19024 6928
rect 10968 6808 11020 6817
rect 12440 6808 12492 6860
rect 17132 6808 17184 6860
rect 21364 6808 21416 6860
rect 22652 6808 22704 6860
rect 24952 6808 25004 6860
rect 8576 6604 8628 6656
rect 8852 6604 8904 6656
rect 9312 6604 9364 6656
rect 9956 6740 10008 6792
rect 12624 6740 12676 6792
rect 11980 6672 12032 6724
rect 11060 6604 11112 6656
rect 12256 6604 12308 6656
rect 13728 6604 13780 6656
rect 14832 6783 14884 6792
rect 14832 6749 14841 6783
rect 14841 6749 14875 6783
rect 14875 6749 14884 6783
rect 14832 6740 14884 6749
rect 15660 6783 15712 6792
rect 15660 6749 15669 6783
rect 15669 6749 15703 6783
rect 15703 6749 15712 6783
rect 15660 6740 15712 6749
rect 17960 6740 18012 6792
rect 18236 6740 18288 6792
rect 19524 6740 19576 6792
rect 24124 6740 24176 6792
rect 25136 6740 25188 6792
rect 21916 6672 21968 6724
rect 14924 6647 14976 6656
rect 14924 6613 14933 6647
rect 14933 6613 14967 6647
rect 14967 6613 14976 6647
rect 14924 6604 14976 6613
rect 15476 6647 15528 6656
rect 15476 6613 15485 6647
rect 15485 6613 15519 6647
rect 15519 6613 15528 6647
rect 15476 6604 15528 6613
rect 17776 6604 17828 6656
rect 22100 6647 22152 6656
rect 22100 6613 22109 6647
rect 22109 6613 22143 6647
rect 22143 6613 22152 6647
rect 22100 6604 22152 6613
rect 25044 6604 25096 6656
rect 8214 6502 8266 6554
rect 8278 6502 8330 6554
rect 8342 6502 8394 6554
rect 8406 6502 8458 6554
rect 8470 6502 8522 6554
rect 16214 6502 16266 6554
rect 16278 6502 16330 6554
rect 16342 6502 16394 6554
rect 16406 6502 16458 6554
rect 16470 6502 16522 6554
rect 24214 6502 24266 6554
rect 24278 6502 24330 6554
rect 24342 6502 24394 6554
rect 24406 6502 24458 6554
rect 24470 6502 24522 6554
rect 1768 6400 1820 6452
rect 3148 6443 3200 6452
rect 3148 6409 3157 6443
rect 3157 6409 3191 6443
rect 3191 6409 3200 6443
rect 3148 6400 3200 6409
rect 4804 6332 4856 6384
rect 4896 6332 4948 6384
rect 3424 6239 3476 6248
rect 3424 6205 3433 6239
rect 3433 6205 3467 6239
rect 3467 6205 3476 6239
rect 3424 6196 3476 6205
rect 3976 6196 4028 6248
rect 5172 6307 5224 6316
rect 5172 6273 5181 6307
rect 5181 6273 5215 6307
rect 5215 6273 5224 6307
rect 5172 6264 5224 6273
rect 5448 6307 5500 6316
rect 5448 6273 5457 6307
rect 5457 6273 5491 6307
rect 5491 6273 5500 6307
rect 5448 6264 5500 6273
rect 6368 6400 6420 6452
rect 7012 6400 7064 6452
rect 5540 6196 5592 6248
rect 7104 6264 7156 6316
rect 10508 6400 10560 6452
rect 11796 6400 11848 6452
rect 12256 6443 12308 6452
rect 12256 6409 12265 6443
rect 12265 6409 12299 6443
rect 12299 6409 12308 6443
rect 12256 6400 12308 6409
rect 7840 6332 7892 6384
rect 8208 6332 8260 6384
rect 8944 6332 8996 6384
rect 9220 6332 9272 6384
rect 9312 6332 9364 6384
rect 8300 6264 8352 6316
rect 8760 6307 8812 6316
rect 8760 6273 8769 6307
rect 8769 6273 8803 6307
rect 8803 6273 8812 6307
rect 8760 6264 8812 6273
rect 8852 6264 8904 6316
rect 9864 6264 9916 6316
rect 9956 6307 10008 6316
rect 9956 6273 9965 6307
rect 9965 6273 9999 6307
rect 9999 6273 10008 6307
rect 9956 6264 10008 6273
rect 11428 6264 11480 6316
rect 12624 6332 12676 6384
rect 13360 6375 13412 6384
rect 13360 6341 13369 6375
rect 13369 6341 13403 6375
rect 13403 6341 13412 6375
rect 13360 6332 13412 6341
rect 13912 6264 13964 6316
rect 15844 6264 15896 6316
rect 16948 6264 17000 6316
rect 17684 6307 17736 6316
rect 17684 6273 17693 6307
rect 17693 6273 17727 6307
rect 17727 6273 17736 6307
rect 17684 6264 17736 6273
rect 8576 6196 8628 6248
rect 10324 6196 10376 6248
rect 2872 6060 2924 6112
rect 7656 6060 7708 6112
rect 7748 6060 7800 6112
rect 8760 6128 8812 6180
rect 9404 6128 9456 6180
rect 9772 6128 9824 6180
rect 13820 6196 13872 6248
rect 14464 6239 14516 6248
rect 14464 6205 14473 6239
rect 14473 6205 14507 6239
rect 14507 6205 14516 6239
rect 14464 6196 14516 6205
rect 15108 6196 15160 6248
rect 18604 6307 18656 6316
rect 18604 6273 18613 6307
rect 18613 6273 18647 6307
rect 18647 6273 18656 6307
rect 18604 6264 18656 6273
rect 19156 6264 19208 6316
rect 21088 6400 21140 6452
rect 21364 6443 21416 6452
rect 21364 6409 21373 6443
rect 21373 6409 21407 6443
rect 21407 6409 21416 6443
rect 21364 6400 21416 6409
rect 25044 6443 25096 6452
rect 25044 6409 25053 6443
rect 25053 6409 25087 6443
rect 25087 6409 25096 6443
rect 25044 6400 25096 6409
rect 22376 6332 22428 6384
rect 23664 6332 23716 6384
rect 22100 6264 22152 6316
rect 19616 6196 19668 6248
rect 20628 6196 20680 6248
rect 20904 6239 20956 6248
rect 20904 6205 20913 6239
rect 20913 6205 20947 6239
rect 20947 6205 20956 6239
rect 20904 6196 20956 6205
rect 23112 6264 23164 6316
rect 22376 6239 22428 6248
rect 22376 6205 22385 6239
rect 22385 6205 22419 6239
rect 22419 6205 22428 6239
rect 22376 6196 22428 6205
rect 22652 6196 22704 6248
rect 23940 6196 23992 6248
rect 8208 6060 8260 6112
rect 8668 6060 8720 6112
rect 9588 6060 9640 6112
rect 10048 6060 10100 6112
rect 15936 6060 15988 6112
rect 17040 6060 17092 6112
rect 17224 6060 17276 6112
rect 18236 6060 18288 6112
rect 19708 6060 19760 6112
rect 19800 6060 19852 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 12214 5958 12266 6010
rect 12278 5958 12330 6010
rect 12342 5958 12394 6010
rect 12406 5958 12458 6010
rect 12470 5958 12522 6010
rect 20214 5958 20266 6010
rect 20278 5958 20330 6010
rect 20342 5958 20394 6010
rect 20406 5958 20458 6010
rect 20470 5958 20522 6010
rect 2780 5831 2832 5840
rect 2780 5797 2789 5831
rect 2789 5797 2823 5831
rect 2823 5797 2832 5831
rect 2780 5788 2832 5797
rect 4712 5788 4764 5840
rect 5172 5856 5224 5908
rect 2504 5652 2556 5704
rect 2872 5652 2924 5704
rect 3332 5695 3384 5704
rect 3332 5661 3371 5695
rect 3371 5661 3384 5695
rect 3332 5652 3384 5661
rect 3516 5695 3568 5704
rect 3516 5661 3518 5695
rect 3518 5661 3552 5695
rect 3552 5661 3568 5695
rect 3516 5652 3568 5661
rect 4712 5695 4764 5704
rect 4712 5661 4721 5695
rect 4721 5661 4755 5695
rect 4755 5661 4764 5695
rect 4712 5652 4764 5661
rect 5172 5652 5224 5704
rect 5264 5695 5316 5704
rect 5264 5661 5273 5695
rect 5273 5661 5307 5695
rect 5307 5661 5316 5695
rect 5264 5652 5316 5661
rect 6092 5652 6144 5704
rect 6920 5788 6972 5840
rect 7104 5899 7156 5908
rect 7104 5865 7113 5899
rect 7113 5865 7147 5899
rect 7147 5865 7156 5899
rect 7104 5856 7156 5865
rect 11428 5856 11480 5908
rect 12072 5856 12124 5908
rect 8944 5788 8996 5840
rect 15108 5899 15160 5908
rect 15108 5865 15117 5899
rect 15117 5865 15151 5899
rect 15151 5865 15160 5899
rect 15108 5856 15160 5865
rect 3240 5584 3292 5636
rect 6000 5584 6052 5636
rect 2044 5559 2096 5568
rect 2044 5525 2053 5559
rect 2053 5525 2087 5559
rect 2087 5525 2096 5559
rect 2044 5516 2096 5525
rect 3148 5559 3200 5568
rect 3148 5525 3157 5559
rect 3157 5525 3191 5559
rect 3191 5525 3200 5559
rect 3148 5516 3200 5525
rect 5908 5516 5960 5568
rect 7012 5584 7064 5636
rect 7104 5627 7156 5636
rect 7104 5593 7113 5627
rect 7113 5593 7147 5627
rect 7147 5593 7156 5627
rect 7104 5584 7156 5593
rect 7380 5695 7432 5704
rect 7380 5661 7389 5695
rect 7389 5661 7423 5695
rect 7423 5661 7432 5695
rect 7380 5652 7432 5661
rect 7840 5652 7892 5704
rect 8300 5720 8352 5772
rect 13636 5788 13688 5840
rect 13728 5788 13780 5840
rect 19432 5856 19484 5908
rect 23664 5899 23716 5908
rect 23664 5865 23673 5899
rect 23673 5865 23707 5899
rect 23707 5865 23716 5899
rect 23664 5856 23716 5865
rect 8208 5695 8260 5704
rect 8208 5661 8217 5695
rect 8217 5661 8251 5695
rect 8251 5661 8260 5695
rect 8208 5652 8260 5661
rect 7564 5584 7616 5636
rect 7656 5516 7708 5568
rect 7748 5516 7800 5568
rect 8024 5584 8076 5636
rect 13268 5720 13320 5772
rect 13820 5720 13872 5772
rect 8760 5652 8812 5704
rect 9036 5695 9088 5704
rect 9036 5661 9045 5695
rect 9045 5661 9079 5695
rect 9079 5661 9088 5695
rect 9036 5652 9088 5661
rect 11428 5652 11480 5704
rect 10048 5584 10100 5636
rect 11980 5584 12032 5636
rect 13360 5627 13412 5636
rect 13360 5593 13369 5627
rect 13369 5593 13403 5627
rect 13403 5593 13412 5627
rect 13360 5584 13412 5593
rect 9496 5516 9548 5568
rect 11520 5559 11572 5568
rect 11520 5525 11529 5559
rect 11529 5525 11563 5559
rect 11563 5525 11572 5559
rect 11520 5516 11572 5525
rect 12072 5516 12124 5568
rect 16120 5763 16172 5772
rect 16120 5729 16129 5763
rect 16129 5729 16163 5763
rect 16163 5729 16172 5763
rect 16120 5720 16172 5729
rect 19524 5763 19576 5772
rect 19524 5729 19533 5763
rect 19533 5729 19567 5763
rect 19567 5729 19576 5763
rect 19524 5720 19576 5729
rect 19800 5763 19852 5772
rect 19800 5729 19809 5763
rect 19809 5729 19843 5763
rect 19843 5729 19852 5763
rect 19800 5720 19852 5729
rect 23388 5695 23440 5704
rect 23388 5661 23397 5695
rect 23397 5661 23431 5695
rect 23431 5661 23440 5695
rect 23388 5652 23440 5661
rect 23572 5652 23624 5704
rect 23756 5652 23808 5704
rect 14464 5584 14516 5636
rect 16672 5584 16724 5636
rect 17224 5627 17276 5636
rect 17224 5593 17233 5627
rect 17233 5593 17267 5627
rect 17267 5593 17276 5627
rect 17224 5584 17276 5593
rect 18236 5584 18288 5636
rect 20812 5584 20864 5636
rect 15936 5559 15988 5568
rect 15936 5525 15945 5559
rect 15945 5525 15979 5559
rect 15979 5525 15988 5559
rect 15936 5516 15988 5525
rect 18144 5516 18196 5568
rect 20168 5516 20220 5568
rect 20628 5516 20680 5568
rect 23296 5516 23348 5568
rect 8214 5414 8266 5466
rect 8278 5414 8330 5466
rect 8342 5414 8394 5466
rect 8406 5414 8458 5466
rect 8470 5414 8522 5466
rect 16214 5414 16266 5466
rect 16278 5414 16330 5466
rect 16342 5414 16394 5466
rect 16406 5414 16458 5466
rect 16470 5414 16522 5466
rect 24214 5414 24266 5466
rect 24278 5414 24330 5466
rect 24342 5414 24394 5466
rect 24406 5414 24458 5466
rect 24470 5414 24522 5466
rect 3240 5312 3292 5364
rect 3608 5312 3660 5364
rect 7012 5312 7064 5364
rect 7656 5312 7708 5364
rect 7840 5312 7892 5364
rect 8944 5312 8996 5364
rect 2044 5244 2096 5296
rect 2780 5244 2832 5296
rect 3792 5244 3844 5296
rect 4804 5287 4856 5296
rect 4804 5253 4813 5287
rect 4813 5253 4847 5287
rect 4847 5253 4856 5287
rect 4804 5244 4856 5253
rect 1492 5219 1544 5228
rect 1492 5185 1501 5219
rect 1501 5185 1535 5219
rect 1535 5185 1544 5219
rect 1492 5176 1544 5185
rect 3332 5176 3384 5228
rect 3516 5108 3568 5160
rect 3976 5108 4028 5160
rect 4528 5219 4580 5228
rect 4528 5185 4537 5219
rect 4537 5185 4571 5219
rect 4571 5185 4580 5219
rect 4528 5176 4580 5185
rect 4712 5219 4764 5228
rect 4712 5185 4719 5219
rect 4719 5185 4764 5219
rect 4712 5176 4764 5185
rect 4896 5219 4948 5228
rect 4896 5185 4905 5219
rect 4905 5185 4939 5219
rect 4939 5185 4948 5219
rect 4896 5176 4948 5185
rect 4988 5219 5040 5228
rect 4988 5185 5021 5219
rect 5021 5185 5040 5219
rect 6000 5219 6052 5228
rect 4988 5176 5040 5185
rect 6000 5185 6008 5219
rect 6008 5185 6042 5219
rect 6042 5185 6052 5219
rect 6000 5176 6052 5185
rect 6920 5244 6972 5296
rect 9128 5244 9180 5296
rect 9588 5287 9640 5296
rect 9588 5253 9597 5287
rect 9597 5253 9631 5287
rect 9631 5253 9640 5287
rect 9588 5244 9640 5253
rect 9864 5312 9916 5364
rect 14924 5312 14976 5364
rect 15752 5355 15804 5364
rect 15752 5321 15761 5355
rect 15761 5321 15795 5355
rect 15795 5321 15804 5355
rect 15752 5312 15804 5321
rect 5080 5040 5132 5092
rect 7564 5219 7616 5228
rect 7564 5185 7573 5219
rect 7573 5185 7607 5219
rect 7607 5185 7616 5219
rect 7564 5176 7616 5185
rect 7932 5176 7984 5228
rect 12624 5244 12676 5296
rect 13360 5244 13412 5296
rect 10324 5219 10376 5228
rect 10324 5185 10333 5219
rect 10333 5185 10367 5219
rect 10367 5185 10376 5219
rect 10324 5176 10376 5185
rect 10968 5176 11020 5228
rect 13728 5176 13780 5228
rect 15476 5244 15528 5296
rect 7380 5108 7432 5160
rect 11888 5151 11940 5160
rect 11888 5117 11897 5151
rect 11897 5117 11931 5151
rect 11931 5117 11940 5151
rect 11888 5108 11940 5117
rect 7104 5040 7156 5092
rect 14188 5040 14240 5092
rect 15108 5219 15160 5228
rect 15108 5185 15117 5219
rect 15117 5185 15151 5219
rect 15151 5185 15160 5219
rect 15108 5176 15160 5185
rect 16120 5312 16172 5364
rect 17684 5312 17736 5364
rect 18144 5312 18196 5364
rect 20168 5312 20220 5364
rect 20812 5312 20864 5364
rect 19708 5244 19760 5296
rect 14924 5108 14976 5160
rect 16028 5219 16080 5228
rect 16028 5185 16036 5219
rect 16036 5185 16070 5219
rect 16070 5185 16080 5219
rect 16028 5176 16080 5185
rect 16120 5219 16172 5228
rect 16120 5185 16129 5219
rect 16129 5185 16163 5219
rect 16163 5185 16172 5219
rect 16120 5176 16172 5185
rect 16948 5176 17000 5228
rect 19156 5219 19208 5228
rect 19156 5185 19165 5219
rect 19165 5185 19199 5219
rect 19199 5185 19208 5219
rect 19156 5176 19208 5185
rect 17040 5108 17092 5160
rect 19984 5176 20036 5228
rect 20628 5176 20680 5228
rect 22376 5312 22428 5364
rect 23664 5244 23716 5296
rect 20076 5108 20128 5160
rect 15200 5040 15252 5092
rect 15844 5040 15896 5092
rect 23112 5219 23164 5228
rect 23112 5185 23121 5219
rect 23121 5185 23155 5219
rect 23155 5185 23164 5219
rect 23112 5176 23164 5185
rect 7012 4972 7064 5024
rect 8484 4972 8536 5024
rect 11980 4972 12032 5024
rect 13820 4972 13872 5024
rect 14556 4972 14608 5024
rect 20720 4972 20772 5024
rect 22652 5108 22704 5160
rect 23112 5040 23164 5092
rect 24952 4972 25004 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 12214 4870 12266 4922
rect 12278 4870 12330 4922
rect 12342 4870 12394 4922
rect 12406 4870 12458 4922
rect 12470 4870 12522 4922
rect 20214 4870 20266 4922
rect 20278 4870 20330 4922
rect 20342 4870 20394 4922
rect 20406 4870 20458 4922
rect 20470 4870 20522 4922
rect 3792 4768 3844 4820
rect 4896 4768 4948 4820
rect 5264 4700 5316 4752
rect 2504 4632 2556 4684
rect 3056 4632 3108 4684
rect 3516 4632 3568 4684
rect 1860 4607 1912 4616
rect 1860 4573 1869 4607
rect 1869 4573 1903 4607
rect 1903 4573 1912 4607
rect 1860 4564 1912 4573
rect 3148 4564 3200 4616
rect 4160 4632 4212 4684
rect 5540 4700 5592 4752
rect 7656 4768 7708 4820
rect 7932 4768 7984 4820
rect 9128 4768 9180 4820
rect 11888 4811 11940 4820
rect 11888 4777 11897 4811
rect 11897 4777 11931 4811
rect 11931 4777 11940 4811
rect 11888 4768 11940 4777
rect 12624 4768 12676 4820
rect 13820 4768 13872 4820
rect 4804 4564 4856 4616
rect 10508 4743 10560 4752
rect 10508 4709 10517 4743
rect 10517 4709 10551 4743
rect 10551 4709 10560 4743
rect 10508 4700 10560 4709
rect 11152 4700 11204 4752
rect 16028 4700 16080 4752
rect 16948 4768 17000 4820
rect 17132 4768 17184 4820
rect 19340 4700 19392 4752
rect 3700 4428 3752 4480
rect 7012 4607 7064 4616
rect 7012 4573 7021 4607
rect 7021 4573 7055 4607
rect 7055 4573 7064 4607
rect 7012 4564 7064 4573
rect 7196 4564 7248 4616
rect 11980 4632 12032 4684
rect 8484 4607 8536 4616
rect 8484 4573 8493 4607
rect 8493 4573 8527 4607
rect 8527 4573 8536 4607
rect 8484 4564 8536 4573
rect 9312 4564 9364 4616
rect 9956 4564 10008 4616
rect 11428 4564 11480 4616
rect 12072 4607 12124 4616
rect 12072 4573 12081 4607
rect 12081 4573 12115 4607
rect 12115 4573 12124 4607
rect 12072 4564 12124 4573
rect 13636 4632 13688 4684
rect 14464 4632 14516 4684
rect 18788 4632 18840 4684
rect 20904 4768 20956 4820
rect 22376 4768 22428 4820
rect 23112 4811 23164 4820
rect 23112 4777 23121 4811
rect 23121 4777 23155 4811
rect 23155 4777 23164 4811
rect 23112 4768 23164 4777
rect 23388 4811 23440 4820
rect 23388 4777 23397 4811
rect 23397 4777 23431 4811
rect 23431 4777 23440 4811
rect 23388 4768 23440 4777
rect 24860 4768 24912 4820
rect 7196 4428 7248 4480
rect 7472 4428 7524 4480
rect 8024 4428 8076 4480
rect 12624 4496 12676 4548
rect 13728 4607 13780 4616
rect 13728 4573 13737 4607
rect 13737 4573 13771 4607
rect 13771 4573 13780 4607
rect 13728 4564 13780 4573
rect 17684 4607 17736 4616
rect 17684 4573 17693 4607
rect 17693 4573 17727 4607
rect 17727 4573 17736 4607
rect 17684 4564 17736 4573
rect 20720 4675 20772 4684
rect 20720 4641 20729 4675
rect 20729 4641 20763 4675
rect 20763 4641 20772 4675
rect 20720 4632 20772 4641
rect 14372 4496 14424 4548
rect 14556 4496 14608 4548
rect 16120 4496 16172 4548
rect 11520 4428 11572 4480
rect 12992 4428 13044 4480
rect 15108 4428 15160 4480
rect 17500 4471 17552 4480
rect 17500 4437 17509 4471
rect 17509 4437 17543 4471
rect 17543 4437 17552 4471
rect 17500 4428 17552 4437
rect 18512 4471 18564 4480
rect 18512 4437 18521 4471
rect 18521 4437 18555 4471
rect 18555 4437 18564 4471
rect 18512 4428 18564 4437
rect 19800 4564 19852 4616
rect 23756 4632 23808 4684
rect 23848 4675 23900 4684
rect 23848 4641 23857 4675
rect 23857 4641 23891 4675
rect 23891 4641 23900 4675
rect 23848 4632 23900 4641
rect 24032 4675 24084 4684
rect 24032 4641 24041 4675
rect 24041 4641 24075 4675
rect 24075 4641 24084 4675
rect 24032 4632 24084 4641
rect 20996 4496 21048 4548
rect 19892 4428 19944 4480
rect 20352 4428 20404 4480
rect 22560 4564 22612 4616
rect 24952 4675 25004 4684
rect 24952 4641 24961 4675
rect 24961 4641 24995 4675
rect 24995 4641 25004 4675
rect 24952 4632 25004 4641
rect 22560 4471 22612 4480
rect 22560 4437 22569 4471
rect 22569 4437 22603 4471
rect 22603 4437 22612 4471
rect 22560 4428 22612 4437
rect 24768 4428 24820 4480
rect 8214 4326 8266 4378
rect 8278 4326 8330 4378
rect 8342 4326 8394 4378
rect 8406 4326 8458 4378
rect 8470 4326 8522 4378
rect 16214 4326 16266 4378
rect 16278 4326 16330 4378
rect 16342 4326 16394 4378
rect 16406 4326 16458 4378
rect 16470 4326 16522 4378
rect 24214 4326 24266 4378
rect 24278 4326 24330 4378
rect 24342 4326 24394 4378
rect 24406 4326 24458 4378
rect 24470 4326 24522 4378
rect 4160 4224 4212 4276
rect 4620 4224 4672 4276
rect 7196 4224 7248 4276
rect 2964 4156 3016 4208
rect 1492 4088 1544 4140
rect 3700 4131 3752 4140
rect 1952 4063 2004 4072
rect 1952 4029 1961 4063
rect 1961 4029 1995 4063
rect 1995 4029 2004 4063
rect 1952 4020 2004 4029
rect 3700 4097 3709 4131
rect 3709 4097 3743 4131
rect 3743 4097 3752 4131
rect 3700 4088 3752 4097
rect 4804 4131 4856 4140
rect 4804 4097 4812 4131
rect 4812 4097 4846 4131
rect 4846 4097 4856 4131
rect 4804 4088 4856 4097
rect 4988 4088 5040 4140
rect 7472 4131 7524 4140
rect 7472 4097 7481 4131
rect 7481 4097 7515 4131
rect 7515 4097 7524 4131
rect 7472 4088 7524 4097
rect 8024 4199 8076 4208
rect 8024 4165 8033 4199
rect 8033 4165 8067 4199
rect 8067 4165 8076 4199
rect 8024 4156 8076 4165
rect 6644 4020 6696 4072
rect 7104 4063 7156 4072
rect 7104 4029 7113 4063
rect 7113 4029 7147 4063
rect 7147 4029 7156 4063
rect 7104 4020 7156 4029
rect 8116 4088 8168 4140
rect 10508 4224 10560 4276
rect 10968 4224 11020 4276
rect 8576 4088 8628 4140
rect 8668 4088 8720 4140
rect 9128 4131 9180 4140
rect 9128 4097 9137 4131
rect 9137 4097 9171 4131
rect 9171 4097 9180 4131
rect 9128 4088 9180 4097
rect 9220 4063 9272 4072
rect 9220 4029 9229 4063
rect 9229 4029 9263 4063
rect 9263 4029 9272 4063
rect 9220 4020 9272 4029
rect 3056 3952 3108 4004
rect 6276 3952 6328 4004
rect 8300 3952 8352 4004
rect 8760 3952 8812 4004
rect 10600 4088 10652 4140
rect 11152 4131 11204 4140
rect 11152 4097 11161 4131
rect 11161 4097 11195 4131
rect 11195 4097 11204 4131
rect 11152 4088 11204 4097
rect 14464 4224 14516 4276
rect 17592 4224 17644 4276
rect 17684 4224 17736 4276
rect 19340 4224 19392 4276
rect 12992 4156 13044 4208
rect 16488 4156 16540 4208
rect 18512 4156 18564 4208
rect 14188 4131 14240 4140
rect 14188 4097 14197 4131
rect 14197 4097 14231 4131
rect 14231 4097 14240 4131
rect 14188 4088 14240 4097
rect 14464 4088 14516 4140
rect 20628 4224 20680 4276
rect 24768 4267 24820 4276
rect 24768 4233 24777 4267
rect 24777 4233 24811 4267
rect 24811 4233 24820 4267
rect 24768 4224 24820 4233
rect 22560 4156 22612 4208
rect 11980 4063 12032 4072
rect 11980 4029 11989 4063
rect 11989 4029 12023 4063
rect 12023 4029 12032 4063
rect 11980 4020 12032 4029
rect 16120 4020 16172 4072
rect 4804 3884 4856 3936
rect 7472 3927 7524 3936
rect 7472 3893 7481 3927
rect 7481 3893 7515 3927
rect 7515 3893 7524 3927
rect 7472 3884 7524 3893
rect 7564 3884 7616 3936
rect 9128 3884 9180 3936
rect 11336 3952 11388 4004
rect 14372 3995 14424 4004
rect 14372 3961 14381 3995
rect 14381 3961 14415 3995
rect 14415 3961 14424 3995
rect 14372 3952 14424 3961
rect 16028 3952 16080 4004
rect 9772 3927 9824 3936
rect 9772 3893 9781 3927
rect 9781 3893 9815 3927
rect 9815 3893 9824 3927
rect 9772 3884 9824 3893
rect 10600 3884 10652 3936
rect 11152 3927 11204 3936
rect 11152 3893 11161 3927
rect 11161 3893 11195 3927
rect 11195 3893 11204 3927
rect 11152 3884 11204 3893
rect 11428 3884 11480 3936
rect 12992 3884 13044 3936
rect 17132 4020 17184 4072
rect 17592 4020 17644 4072
rect 20352 4131 20404 4140
rect 20352 4097 20361 4131
rect 20361 4097 20395 4131
rect 20395 4097 20404 4131
rect 20352 4088 20404 4097
rect 20812 4131 20864 4140
rect 20812 4097 20821 4131
rect 20821 4097 20855 4131
rect 20855 4097 20864 4131
rect 20812 4088 20864 4097
rect 16672 3952 16724 4004
rect 18052 3884 18104 3936
rect 19616 3952 19668 4004
rect 23020 4131 23072 4140
rect 23020 4097 23029 4131
rect 23029 4097 23063 4131
rect 23063 4097 23072 4131
rect 23020 4088 23072 4097
rect 23296 4063 23348 4072
rect 23296 4029 23305 4063
rect 23305 4029 23339 4063
rect 23339 4029 23348 4063
rect 23296 4020 23348 4029
rect 20996 3995 21048 4004
rect 20996 3961 21005 3995
rect 21005 3961 21039 3995
rect 21039 3961 21048 3995
rect 20996 3952 21048 3961
rect 19800 3884 19852 3936
rect 19892 3927 19944 3936
rect 19892 3893 19901 3927
rect 19901 3893 19935 3927
rect 19935 3893 19944 3927
rect 19892 3884 19944 3893
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 12214 3782 12266 3834
rect 12278 3782 12330 3834
rect 12342 3782 12394 3834
rect 12406 3782 12458 3834
rect 12470 3782 12522 3834
rect 20214 3782 20266 3834
rect 20278 3782 20330 3834
rect 20342 3782 20394 3834
rect 20406 3782 20458 3834
rect 20470 3782 20522 3834
rect 1952 3680 2004 3732
rect 2964 3680 3016 3732
rect 6644 3723 6696 3732
rect 6644 3689 6653 3723
rect 6653 3689 6687 3723
rect 6687 3689 6696 3723
rect 6644 3680 6696 3689
rect 7380 3723 7432 3732
rect 7380 3689 7389 3723
rect 7389 3689 7423 3723
rect 7423 3689 7432 3723
rect 7380 3680 7432 3689
rect 6184 3612 6236 3664
rect 7472 3612 7524 3664
rect 4804 3544 4856 3596
rect 2872 3476 2924 3528
rect 2504 3408 2556 3460
rect 6184 3519 6236 3528
rect 6184 3485 6192 3519
rect 6192 3485 6226 3519
rect 6226 3485 6236 3519
rect 6184 3476 6236 3485
rect 6276 3519 6328 3528
rect 6276 3485 6285 3519
rect 6285 3485 6319 3519
rect 6319 3485 6328 3519
rect 6276 3476 6328 3485
rect 7564 3519 7616 3528
rect 7564 3485 7573 3519
rect 7573 3485 7607 3519
rect 7607 3485 7616 3519
rect 7564 3476 7616 3485
rect 7748 3519 7800 3528
rect 7748 3485 7757 3519
rect 7757 3485 7791 3519
rect 7791 3485 7800 3519
rect 7748 3476 7800 3485
rect 8852 3680 8904 3732
rect 10508 3680 10560 3732
rect 11336 3680 11388 3732
rect 11980 3680 12032 3732
rect 16488 3723 16540 3732
rect 16488 3689 16497 3723
rect 16497 3689 16531 3723
rect 16531 3689 16540 3723
rect 16488 3680 16540 3689
rect 17592 3680 17644 3732
rect 20628 3680 20680 3732
rect 8300 3519 8352 3528
rect 8300 3485 8309 3519
rect 8309 3485 8343 3519
rect 8343 3485 8352 3519
rect 8300 3476 8352 3485
rect 9036 3544 9088 3596
rect 9864 3544 9916 3596
rect 10968 3544 11020 3596
rect 10600 3476 10652 3528
rect 13084 3612 13136 3664
rect 13268 3587 13320 3596
rect 13268 3553 13277 3587
rect 13277 3553 13311 3587
rect 13311 3553 13320 3587
rect 13268 3544 13320 3553
rect 12992 3476 13044 3528
rect 2872 3340 2924 3392
rect 3608 3340 3660 3392
rect 9220 3408 9272 3460
rect 9772 3408 9824 3460
rect 12072 3408 12124 3460
rect 14556 3476 14608 3528
rect 15936 3544 15988 3596
rect 16672 3612 16724 3664
rect 21088 3612 21140 3664
rect 17500 3587 17552 3596
rect 17500 3553 17509 3587
rect 17509 3553 17543 3587
rect 17543 3553 17552 3587
rect 17500 3544 17552 3553
rect 18052 3544 18104 3596
rect 23020 3544 23072 3596
rect 4620 3340 4672 3392
rect 9312 3340 9364 3392
rect 14188 3340 14240 3392
rect 15016 3340 15068 3392
rect 16672 3519 16724 3528
rect 16672 3485 16681 3519
rect 16681 3485 16715 3519
rect 16715 3485 16724 3519
rect 16672 3476 16724 3485
rect 19340 3519 19392 3528
rect 19340 3485 19349 3519
rect 19349 3485 19383 3519
rect 19383 3485 19392 3519
rect 19340 3476 19392 3485
rect 20076 3476 20128 3528
rect 23664 3680 23716 3732
rect 23572 3519 23624 3528
rect 19708 3408 19760 3460
rect 20628 3408 20680 3460
rect 23572 3485 23581 3519
rect 23581 3485 23615 3519
rect 23615 3485 23624 3519
rect 23572 3476 23624 3485
rect 23756 3519 23808 3528
rect 23756 3485 23765 3519
rect 23765 3485 23799 3519
rect 23799 3485 23808 3519
rect 23756 3476 23808 3485
rect 22008 3408 22060 3460
rect 21456 3340 21508 3392
rect 21548 3340 21600 3392
rect 8214 3238 8266 3290
rect 8278 3238 8330 3290
rect 8342 3238 8394 3290
rect 8406 3238 8458 3290
rect 8470 3238 8522 3290
rect 16214 3238 16266 3290
rect 16278 3238 16330 3290
rect 16342 3238 16394 3290
rect 16406 3238 16458 3290
rect 16470 3238 16522 3290
rect 24214 3238 24266 3290
rect 24278 3238 24330 3290
rect 24342 3238 24394 3290
rect 24406 3238 24458 3290
rect 24470 3238 24522 3290
rect 4712 3136 4764 3188
rect 5172 3136 5224 3188
rect 2504 3000 2556 3052
rect 3608 3043 3660 3052
rect 3608 3009 3617 3043
rect 3617 3009 3651 3043
rect 3651 3009 3660 3043
rect 3608 3000 3660 3009
rect 4804 2932 4856 2984
rect 4988 2975 5040 2984
rect 4988 2941 4997 2975
rect 4997 2941 5031 2975
rect 5031 2941 5040 2975
rect 4988 2932 5040 2941
rect 5632 2932 5684 2984
rect 4068 2864 4120 2916
rect 1492 2796 1544 2848
rect 2872 2796 2924 2848
rect 3976 2796 4028 2848
rect 8116 3136 8168 3188
rect 9496 3136 9548 3188
rect 14188 3136 14240 3188
rect 16212 3136 16264 3188
rect 5908 3043 5960 3052
rect 5908 3009 5917 3043
rect 5917 3009 5951 3043
rect 5951 3009 5960 3043
rect 5908 3000 5960 3009
rect 6736 3068 6788 3120
rect 7564 3000 7616 3052
rect 9312 3111 9364 3120
rect 9312 3077 9321 3111
rect 9321 3077 9355 3111
rect 9355 3077 9364 3111
rect 9312 3068 9364 3077
rect 11152 3068 11204 3120
rect 6000 2932 6052 2984
rect 7196 2864 7248 2916
rect 7380 2932 7432 2984
rect 9036 3043 9088 3052
rect 9036 3009 9045 3043
rect 9045 3009 9079 3043
rect 9079 3009 9088 3043
rect 9036 3000 9088 3009
rect 9404 2932 9456 2984
rect 12624 3043 12676 3052
rect 12624 3009 12633 3043
rect 12633 3009 12667 3043
rect 12667 3009 12676 3043
rect 12624 3000 12676 3009
rect 12900 3000 12952 3052
rect 13084 3000 13136 3052
rect 14648 3068 14700 3120
rect 17592 3136 17644 3188
rect 21548 3179 21600 3188
rect 21548 3145 21557 3179
rect 21557 3145 21591 3179
rect 21591 3145 21600 3179
rect 21548 3136 21600 3145
rect 22008 3179 22060 3188
rect 22008 3145 22017 3179
rect 22017 3145 22051 3179
rect 22051 3145 22060 3179
rect 22008 3136 22060 3145
rect 13820 3000 13872 3052
rect 14280 3000 14332 3052
rect 12072 2864 12124 2916
rect 15660 3000 15712 3052
rect 7288 2839 7340 2848
rect 7288 2805 7297 2839
rect 7297 2805 7331 2839
rect 7331 2805 7340 2839
rect 7288 2796 7340 2805
rect 9312 2796 9364 2848
rect 11244 2796 11296 2848
rect 12808 2839 12860 2848
rect 12808 2805 12817 2839
rect 12817 2805 12851 2839
rect 12851 2805 12860 2839
rect 12808 2796 12860 2805
rect 14372 2839 14424 2848
rect 14372 2805 14381 2839
rect 14381 2805 14415 2839
rect 14415 2805 14424 2839
rect 14372 2796 14424 2805
rect 14648 2839 14700 2848
rect 14648 2805 14657 2839
rect 14657 2805 14691 2839
rect 14691 2805 14700 2839
rect 14648 2796 14700 2805
rect 14924 2796 14976 2848
rect 21088 3068 21140 3120
rect 15844 3000 15896 3052
rect 16672 3000 16724 3052
rect 19708 3000 19760 3052
rect 19800 3043 19852 3052
rect 19800 3009 19809 3043
rect 19809 3009 19843 3043
rect 19843 3009 19852 3043
rect 19800 3000 19852 3009
rect 21456 3000 21508 3052
rect 23756 3000 23808 3052
rect 16948 2932 17000 2984
rect 16580 2796 16632 2848
rect 17040 2864 17092 2916
rect 17224 2932 17276 2984
rect 19616 2932 19668 2984
rect 20076 2975 20128 2984
rect 20076 2941 20085 2975
rect 20085 2941 20119 2975
rect 20119 2941 20128 2975
rect 20076 2932 20128 2941
rect 18512 2864 18564 2916
rect 18420 2796 18472 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 12214 2694 12266 2746
rect 12278 2694 12330 2746
rect 12342 2694 12394 2746
rect 12406 2694 12458 2746
rect 12470 2694 12522 2746
rect 20214 2694 20266 2746
rect 20278 2694 20330 2746
rect 20342 2694 20394 2746
rect 20406 2694 20458 2746
rect 20470 2694 20522 2746
rect 8576 2592 8628 2644
rect 12624 2592 12676 2644
rect 2872 2456 2924 2508
rect 7012 2499 7064 2508
rect 7012 2465 7021 2499
rect 7021 2465 7055 2499
rect 7055 2465 7064 2499
rect 7012 2456 7064 2465
rect 7196 2456 7248 2508
rect 3148 2252 3200 2304
rect 6000 2388 6052 2440
rect 7472 2388 7524 2440
rect 9864 2456 9916 2508
rect 10876 2499 10928 2508
rect 10876 2465 10885 2499
rect 10885 2465 10919 2499
rect 10919 2465 10928 2499
rect 10876 2456 10928 2465
rect 4436 2320 4488 2372
rect 4620 2320 4672 2372
rect 6276 2252 6328 2304
rect 6460 2320 6512 2372
rect 6736 2363 6788 2372
rect 6736 2329 6745 2363
rect 6745 2329 6779 2363
rect 6779 2329 6788 2363
rect 6736 2320 6788 2329
rect 9128 2388 9180 2440
rect 13084 2388 13136 2440
rect 13728 2592 13780 2644
rect 14188 2635 14240 2644
rect 14188 2601 14197 2635
rect 14197 2601 14231 2635
rect 14231 2601 14240 2635
rect 14188 2592 14240 2601
rect 16212 2635 16264 2644
rect 16212 2601 16221 2635
rect 16221 2601 16255 2635
rect 16255 2601 16264 2635
rect 16212 2592 16264 2601
rect 13728 2388 13780 2440
rect 13912 2456 13964 2508
rect 14280 2456 14332 2508
rect 15660 2499 15712 2508
rect 15660 2465 15669 2499
rect 15669 2465 15703 2499
rect 15703 2465 15712 2499
rect 15660 2456 15712 2465
rect 15936 2499 15988 2508
rect 15936 2465 15945 2499
rect 15945 2465 15979 2499
rect 15979 2465 15988 2499
rect 15936 2456 15988 2465
rect 16672 2456 16724 2508
rect 19892 2456 19944 2508
rect 19984 2499 20036 2508
rect 19984 2465 19993 2499
rect 19993 2465 20027 2499
rect 20027 2465 20036 2499
rect 19984 2456 20036 2465
rect 16580 2388 16632 2440
rect 11152 2363 11204 2372
rect 11152 2329 11161 2363
rect 11161 2329 11195 2363
rect 11195 2329 11204 2363
rect 11152 2320 11204 2329
rect 12808 2320 12860 2372
rect 6828 2295 6880 2304
rect 6828 2261 6837 2295
rect 6837 2261 6871 2295
rect 6871 2261 6880 2295
rect 6828 2252 6880 2261
rect 8116 2295 8168 2304
rect 8116 2261 8125 2295
rect 8125 2261 8159 2295
rect 8159 2261 8168 2295
rect 8116 2252 8168 2261
rect 12164 2252 12216 2304
rect 17500 2252 17552 2304
rect 17776 2320 17828 2372
rect 18420 2431 18472 2440
rect 18420 2397 18429 2431
rect 18429 2397 18463 2431
rect 18463 2397 18472 2431
rect 18420 2388 18472 2397
rect 19064 2252 19116 2304
rect 19616 2388 19668 2440
rect 20628 2388 20680 2440
rect 19708 2295 19760 2304
rect 19708 2261 19717 2295
rect 19717 2261 19751 2295
rect 19751 2261 19760 2295
rect 19708 2252 19760 2261
rect 20444 2295 20496 2304
rect 20444 2261 20453 2295
rect 20453 2261 20487 2295
rect 20487 2261 20496 2295
rect 20444 2252 20496 2261
rect 8214 2150 8266 2202
rect 8278 2150 8330 2202
rect 8342 2150 8394 2202
rect 8406 2150 8458 2202
rect 8470 2150 8522 2202
rect 16214 2150 16266 2202
rect 16278 2150 16330 2202
rect 16342 2150 16394 2202
rect 16406 2150 16458 2202
rect 16470 2150 16522 2202
rect 24214 2150 24266 2202
rect 24278 2150 24330 2202
rect 24342 2150 24394 2202
rect 24406 2150 24458 2202
rect 24470 2150 24522 2202
rect 4896 2091 4948 2100
rect 4896 2057 4905 2091
rect 4905 2057 4939 2091
rect 4939 2057 4948 2091
rect 4896 2048 4948 2057
rect 5632 2091 5684 2100
rect 5632 2057 5641 2091
rect 5641 2057 5675 2091
rect 5675 2057 5684 2091
rect 5632 2048 5684 2057
rect 7748 2048 7800 2100
rect 9496 2091 9548 2100
rect 9496 2057 9505 2091
rect 9505 2057 9539 2091
rect 9539 2057 9548 2091
rect 9496 2048 9548 2057
rect 3148 2023 3200 2032
rect 3148 1989 3157 2023
rect 3157 1989 3191 2023
rect 3191 1989 3200 2023
rect 3148 1980 3200 1989
rect 4160 1980 4212 2032
rect 4436 1980 4488 2032
rect 2872 1955 2924 1964
rect 2872 1921 2881 1955
rect 2881 1921 2915 1955
rect 2915 1921 2924 1955
rect 2872 1912 2924 1921
rect 5908 1955 5960 1964
rect 5908 1921 5916 1955
rect 5916 1921 5950 1955
rect 5950 1921 5960 1955
rect 5908 1912 5960 1921
rect 6000 1955 6052 1964
rect 6000 1921 6009 1955
rect 6009 1921 6043 1955
rect 6043 1921 6052 1955
rect 10876 1980 10928 2032
rect 12164 2048 12216 2100
rect 16672 2048 16724 2100
rect 6000 1912 6052 1921
rect 7288 1912 7340 1964
rect 7564 1955 7616 1964
rect 7564 1921 7573 1955
rect 7573 1921 7607 1955
rect 7607 1921 7616 1955
rect 7564 1912 7616 1921
rect 8668 1955 8720 1964
rect 8668 1921 8677 1955
rect 8677 1921 8711 1955
rect 8711 1921 8720 1955
rect 8668 1912 8720 1921
rect 14372 1980 14424 2032
rect 15016 2023 15068 2032
rect 15016 1989 15025 2023
rect 15025 1989 15059 2023
rect 15059 1989 15068 2023
rect 15016 1980 15068 1989
rect 12072 1912 12124 1964
rect 12900 1955 12952 1964
rect 12900 1921 12909 1955
rect 12909 1921 12943 1955
rect 12943 1921 12952 1955
rect 12900 1912 12952 1921
rect 13084 1955 13136 1964
rect 13084 1921 13093 1955
rect 13093 1921 13127 1955
rect 13127 1921 13136 1955
rect 13084 1912 13136 1921
rect 17776 2048 17828 2100
rect 18512 2091 18564 2100
rect 18512 2057 18521 2091
rect 18521 2057 18555 2091
rect 18555 2057 18564 2091
rect 18512 2048 18564 2057
rect 17500 1980 17552 2032
rect 19064 2023 19116 2032
rect 19064 1989 19073 2023
rect 19073 1989 19107 2023
rect 19107 1989 19116 2023
rect 19064 1980 19116 1989
rect 20444 1980 20496 2032
rect 4896 1844 4948 1896
rect 5080 1819 5132 1828
rect 5080 1785 5089 1819
rect 5089 1785 5123 1819
rect 5123 1785 5132 1819
rect 5080 1776 5132 1785
rect 6276 1844 6328 1896
rect 6736 1844 6788 1896
rect 6460 1776 6512 1828
rect 7380 1887 7432 1896
rect 7380 1853 7389 1887
rect 7389 1853 7423 1887
rect 7423 1853 7432 1887
rect 7380 1844 7432 1853
rect 7472 1887 7524 1896
rect 7472 1853 7481 1887
rect 7481 1853 7515 1887
rect 7515 1853 7524 1887
rect 7472 1844 7524 1853
rect 8392 1844 8444 1896
rect 9220 1844 9272 1896
rect 10968 1887 11020 1896
rect 10968 1853 10977 1887
rect 10977 1853 11011 1887
rect 11011 1853 11020 1887
rect 10968 1844 11020 1853
rect 17040 1887 17092 1896
rect 17040 1853 17049 1887
rect 17049 1853 17083 1887
rect 17083 1853 17092 1887
rect 17040 1844 17092 1853
rect 17776 1844 17828 1896
rect 8852 1708 8904 1760
rect 11796 1708 11848 1760
rect 13544 1751 13596 1760
rect 13544 1717 13553 1751
rect 13553 1717 13587 1751
rect 13587 1717 13596 1751
rect 13544 1708 13596 1717
rect 19708 1708 19760 1760
rect 4214 1606 4266 1658
rect 4278 1606 4330 1658
rect 4342 1606 4394 1658
rect 4406 1606 4458 1658
rect 4470 1606 4522 1658
rect 12214 1606 12266 1658
rect 12278 1606 12330 1658
rect 12342 1606 12394 1658
rect 12406 1606 12458 1658
rect 12470 1606 12522 1658
rect 20214 1606 20266 1658
rect 20278 1606 20330 1658
rect 20342 1606 20394 1658
rect 20406 1606 20458 1658
rect 20470 1606 20522 1658
rect 4988 1504 5040 1556
rect 6828 1547 6880 1556
rect 6828 1513 6837 1547
rect 6837 1513 6871 1547
rect 6871 1513 6880 1547
rect 6828 1504 6880 1513
rect 8392 1547 8444 1556
rect 8392 1513 8401 1547
rect 8401 1513 8435 1547
rect 8435 1513 8444 1547
rect 8392 1504 8444 1513
rect 10968 1504 11020 1556
rect 11152 1504 11204 1556
rect 17040 1547 17092 1556
rect 17040 1513 17049 1547
rect 17049 1513 17083 1547
rect 17083 1513 17092 1547
rect 17040 1504 17092 1513
rect 8668 1436 8720 1488
rect 12072 1436 12124 1488
rect 14924 1436 14976 1488
rect 848 1368 900 1420
rect 7380 1368 7432 1420
rect 8116 1368 8168 1420
rect 2872 1300 2924 1352
rect 4896 1343 4948 1352
rect 4896 1309 4904 1343
rect 4904 1309 4938 1343
rect 4938 1309 4948 1343
rect 4896 1300 4948 1309
rect 5080 1300 5132 1352
rect 6736 1300 6788 1352
rect 9220 1300 9272 1352
rect 11244 1343 11296 1352
rect 11244 1309 11253 1343
rect 11253 1309 11287 1343
rect 11287 1309 11296 1343
rect 11244 1300 11296 1309
rect 11796 1343 11848 1352
rect 11796 1309 11805 1343
rect 11805 1309 11839 1343
rect 11839 1309 11848 1343
rect 11796 1300 11848 1309
rect 13544 1300 13596 1352
rect 15108 1232 15160 1284
rect 14556 1207 14608 1216
rect 14556 1173 14565 1207
rect 14565 1173 14599 1207
rect 14599 1173 14608 1207
rect 14556 1164 14608 1173
rect 18512 1300 18564 1352
rect 19708 1368 19760 1420
rect 8214 1062 8266 1114
rect 8278 1062 8330 1114
rect 8342 1062 8394 1114
rect 8406 1062 8458 1114
rect 8470 1062 8522 1114
rect 16214 1062 16266 1114
rect 16278 1062 16330 1114
rect 16342 1062 16394 1114
rect 16406 1062 16458 1114
rect 16470 1062 16522 1114
rect 24214 1062 24266 1114
rect 24278 1062 24330 1114
rect 24342 1062 24394 1114
rect 24406 1062 24458 1114
rect 24470 1062 24522 1114
<< metal2 >>
rect 1306 21298 1362 22000
rect 1400 21344 1452 21350
rect 1306 21292 1400 21298
rect 1306 21286 1452 21292
rect 3330 21298 3386 22000
rect 1306 21270 1440 21286
rect 3330 21282 3648 21298
rect 3330 21276 3660 21282
rect 3330 21270 3608 21276
rect 1306 21200 1362 21270
rect 3330 21200 3386 21270
rect 3608 21218 3660 21224
rect 5354 21208 5410 22000
rect 5354 21200 5356 21208
rect 5408 21200 5410 21208
rect 7378 21200 7434 22000
rect 9402 21200 9458 22000
rect 11426 21200 11482 22000
rect 13176 21344 13228 21350
rect 13176 21286 13228 21292
rect 5356 21150 5408 21156
rect 7392 20942 7420 21200
rect 9128 21004 9180 21010
rect 9128 20946 9180 20952
rect 7380 20936 7432 20942
rect 7380 20878 7432 20884
rect 6734 20768 6790 20777
rect 6734 20703 6790 20712
rect 4712 20460 4764 20466
rect 4712 20402 4764 20408
rect 4896 20460 4948 20466
rect 4896 20402 4948 20408
rect 204 20392 256 20398
rect 204 20334 256 20340
rect 216 2553 244 20334
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4618 19680 4674 19689
rect 4618 19615 4674 19624
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 3240 18760 3292 18766
rect 3240 18702 3292 18708
rect 4528 18760 4580 18766
rect 4528 18702 4580 18708
rect 3252 18426 3280 18702
rect 4068 18692 4120 18698
rect 4068 18634 4120 18640
rect 3974 18592 4030 18601
rect 3974 18527 4030 18536
rect 3240 18420 3292 18426
rect 3240 18362 3292 18368
rect 3884 17128 3936 17134
rect 3884 17070 3936 17076
rect 3896 16794 3924 17070
rect 3884 16788 3936 16794
rect 3884 16730 3936 16736
rect 3988 16590 4016 18527
rect 4080 18426 4108 18634
rect 4436 18624 4488 18630
rect 4436 18566 4488 18572
rect 4068 18420 4120 18426
rect 4068 18362 4120 18368
rect 4448 18358 4476 18566
rect 4436 18352 4488 18358
rect 4436 18294 4488 18300
rect 4252 18284 4304 18290
rect 4252 18226 4304 18232
rect 4264 18086 4292 18226
rect 4540 18222 4568 18702
rect 4632 18426 4660 19615
rect 4724 19446 4752 20402
rect 4908 19854 4936 20402
rect 5172 20392 5224 20398
rect 5172 20334 5224 20340
rect 4896 19848 4948 19854
rect 4896 19790 4948 19796
rect 4712 19440 4764 19446
rect 4712 19382 4764 19388
rect 4804 19372 4856 19378
rect 4804 19314 4856 19320
rect 4816 18970 4844 19314
rect 4908 18970 4936 19790
rect 5184 19242 5212 20334
rect 5356 20256 5408 20262
rect 5356 20198 5408 20204
rect 5540 20256 5592 20262
rect 5540 20198 5592 20204
rect 5908 20256 5960 20262
rect 5908 20198 5960 20204
rect 5368 19514 5396 20198
rect 5448 19848 5500 19854
rect 5448 19790 5500 19796
rect 5460 19514 5488 19790
rect 5356 19508 5408 19514
rect 5356 19450 5408 19456
rect 5448 19508 5500 19514
rect 5448 19450 5500 19456
rect 5552 19310 5580 20198
rect 5920 19922 5948 20198
rect 5908 19916 5960 19922
rect 5908 19858 5960 19864
rect 5816 19372 5868 19378
rect 5816 19314 5868 19320
rect 5540 19304 5592 19310
rect 5540 19246 5592 19252
rect 5172 19236 5224 19242
rect 5172 19178 5224 19184
rect 5828 18970 5856 19314
rect 4804 18964 4856 18970
rect 4804 18906 4856 18912
rect 4896 18964 4948 18970
rect 4896 18906 4948 18912
rect 5816 18964 5868 18970
rect 5816 18906 5868 18912
rect 5724 18760 5776 18766
rect 5724 18702 5776 18708
rect 6552 18760 6604 18766
rect 6552 18702 6604 18708
rect 5736 18426 5764 18702
rect 5816 18624 5868 18630
rect 5816 18566 5868 18572
rect 6460 18624 6512 18630
rect 6460 18566 6512 18572
rect 4620 18420 4672 18426
rect 4620 18362 4672 18368
rect 4712 18420 4764 18426
rect 4712 18362 4764 18368
rect 5724 18420 5776 18426
rect 5724 18362 5776 18368
rect 4528 18216 4580 18222
rect 4528 18158 4580 18164
rect 4724 18154 4752 18362
rect 5080 18216 5132 18222
rect 5080 18158 5132 18164
rect 4712 18148 4764 18154
rect 4712 18090 4764 18096
rect 4068 18080 4120 18086
rect 4068 18022 4120 18028
rect 4252 18080 4304 18086
rect 4252 18022 4304 18028
rect 4080 17796 4108 18022
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4988 17876 5040 17882
rect 4988 17818 5040 17824
rect 4344 17808 4396 17814
rect 4080 17768 4344 17796
rect 4344 17750 4396 17756
rect 4436 17672 4488 17678
rect 4712 17672 4764 17678
rect 4488 17632 4568 17660
rect 4436 17614 4488 17620
rect 4344 17604 4396 17610
rect 4344 17546 4396 17552
rect 4356 17270 4384 17546
rect 4436 17536 4488 17542
rect 4436 17478 4488 17484
rect 4448 17270 4476 17478
rect 4540 17270 4568 17632
rect 4712 17614 4764 17620
rect 4724 17338 4752 17614
rect 4712 17332 4764 17338
rect 4712 17274 4764 17280
rect 4344 17264 4396 17270
rect 4344 17206 4396 17212
rect 4436 17264 4488 17270
rect 4436 17206 4488 17212
rect 4528 17264 4580 17270
rect 4528 17206 4580 17212
rect 5000 17202 5028 17818
rect 5092 17814 5120 18158
rect 5828 18154 5856 18566
rect 5816 18148 5868 18154
rect 5816 18090 5868 18096
rect 5356 18080 5408 18086
rect 5356 18022 5408 18028
rect 5368 17882 5396 18022
rect 5356 17876 5408 17882
rect 5356 17818 5408 17824
rect 5080 17808 5132 17814
rect 5080 17750 5132 17756
rect 5828 17678 5856 18090
rect 5632 17672 5684 17678
rect 5816 17672 5868 17678
rect 5632 17614 5684 17620
rect 5736 17632 5816 17660
rect 5644 17513 5672 17614
rect 5630 17504 5686 17513
rect 5630 17439 5686 17448
rect 4988 17196 5040 17202
rect 4988 17138 5040 17144
rect 4712 17128 4764 17134
rect 4712 17070 4764 17076
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4724 16794 4752 17070
rect 4712 16788 4764 16794
rect 4712 16730 4764 16736
rect 5000 16590 5028 17138
rect 3976 16584 4028 16590
rect 3976 16526 4028 16532
rect 4252 16584 4304 16590
rect 4252 16526 4304 16532
rect 4988 16584 5040 16590
rect 4988 16526 5040 16532
rect 4160 16448 4212 16454
rect 4160 16390 4212 16396
rect 4172 16114 4200 16390
rect 4264 16182 4292 16526
rect 5736 16454 5764 17632
rect 5816 17614 5868 17620
rect 5816 17536 5868 17542
rect 5816 17478 5868 17484
rect 6184 17536 6236 17542
rect 6184 17478 6236 17484
rect 5828 17202 5856 17478
rect 5816 17196 5868 17202
rect 5816 17138 5868 17144
rect 6092 17196 6144 17202
rect 6196 17184 6224 17478
rect 6144 17156 6224 17184
rect 6092 17138 6144 17144
rect 5828 16590 5856 17138
rect 5908 16992 5960 16998
rect 5908 16934 5960 16940
rect 5920 16726 5948 16934
rect 5908 16720 5960 16726
rect 5908 16662 5960 16668
rect 5816 16584 5868 16590
rect 5816 16526 5868 16532
rect 5724 16448 5776 16454
rect 5724 16390 5776 16396
rect 4252 16176 4304 16182
rect 4252 16118 4304 16124
rect 3424 16108 3476 16114
rect 3424 16050 3476 16056
rect 4160 16108 4212 16114
rect 4160 16050 4212 16056
rect 3056 16040 3108 16046
rect 3056 15982 3108 15988
rect 3068 15638 3096 15982
rect 3148 15904 3200 15910
rect 3148 15846 3200 15852
rect 3056 15632 3108 15638
rect 3056 15574 3108 15580
rect 3056 15496 3108 15502
rect 3056 15438 3108 15444
rect 2964 15360 3016 15366
rect 2964 15302 3016 15308
rect 2976 15094 3004 15302
rect 2964 15088 3016 15094
rect 2964 15030 3016 15036
rect 1492 14952 1544 14958
rect 1492 14894 1544 14900
rect 2688 14952 2740 14958
rect 2688 14894 2740 14900
rect 1504 14414 1532 14894
rect 2136 14476 2188 14482
rect 2136 14418 2188 14424
rect 1492 14408 1544 14414
rect 1492 14350 1544 14356
rect 1504 11694 1532 14350
rect 2148 13938 2176 14418
rect 2136 13932 2188 13938
rect 2136 13874 2188 13880
rect 2700 13870 2728 14894
rect 3068 14550 3096 15438
rect 3056 14544 3108 14550
rect 3056 14486 3108 14492
rect 2964 14272 3016 14278
rect 2964 14214 3016 14220
rect 2688 13864 2740 13870
rect 2688 13806 2740 13812
rect 2976 13530 3004 14214
rect 3068 14074 3096 14486
rect 3160 14414 3188 15846
rect 3436 15706 3464 16050
rect 4620 15904 4672 15910
rect 4620 15846 4672 15852
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 3424 15700 3476 15706
rect 3424 15642 3476 15648
rect 3240 15564 3292 15570
rect 3240 15506 3292 15512
rect 3252 15094 3280 15506
rect 3884 15496 3936 15502
rect 3884 15438 3936 15444
rect 3896 15162 3924 15438
rect 4632 15434 4660 15846
rect 5736 15638 5764 16390
rect 6104 16114 6132 17138
rect 6276 16516 6328 16522
rect 6276 16458 6328 16464
rect 6092 16108 6144 16114
rect 6092 16050 6144 16056
rect 6092 15904 6144 15910
rect 6092 15846 6144 15852
rect 5724 15632 5776 15638
rect 5724 15574 5776 15580
rect 6104 15502 6132 15846
rect 6288 15706 6316 16458
rect 6276 15700 6328 15706
rect 6276 15642 6328 15648
rect 6092 15496 6144 15502
rect 6092 15438 6144 15444
rect 4620 15428 4672 15434
rect 4620 15370 4672 15376
rect 4988 15360 5040 15366
rect 4988 15302 5040 15308
rect 3884 15156 3936 15162
rect 3884 15098 3936 15104
rect 3240 15088 3292 15094
rect 4068 15088 4120 15094
rect 3292 15036 3372 15042
rect 3240 15030 3372 15036
rect 4068 15030 4120 15036
rect 3252 15014 3372 15030
rect 3240 14952 3292 14958
rect 3240 14894 3292 14900
rect 3148 14408 3200 14414
rect 3148 14350 3200 14356
rect 3056 14068 3108 14074
rect 3056 14010 3108 14016
rect 2964 13524 3016 13530
rect 2964 13466 3016 13472
rect 3252 13326 3280 14894
rect 3344 13802 3372 15014
rect 3976 15020 4028 15026
rect 3976 14962 4028 14968
rect 3424 14816 3476 14822
rect 3424 14758 3476 14764
rect 3516 14816 3568 14822
rect 3516 14758 3568 14764
rect 3436 13870 3464 14758
rect 3528 14006 3556 14758
rect 3608 14272 3660 14278
rect 3608 14214 3660 14220
rect 3884 14272 3936 14278
rect 3884 14214 3936 14220
rect 3620 14006 3648 14214
rect 3896 14074 3924 14214
rect 3884 14068 3936 14074
rect 3884 14010 3936 14016
rect 3516 14000 3568 14006
rect 3516 13942 3568 13948
rect 3608 14000 3660 14006
rect 3608 13942 3660 13948
rect 3424 13864 3476 13870
rect 3424 13806 3476 13812
rect 3332 13796 3384 13802
rect 3332 13738 3384 13744
rect 3344 13394 3372 13738
rect 3332 13388 3384 13394
rect 3332 13330 3384 13336
rect 3620 13326 3648 13942
rect 3988 13734 4016 14962
rect 4080 14618 4108 15030
rect 4804 15020 4856 15026
rect 4804 14962 4856 14968
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4068 14612 4120 14618
rect 4068 14554 4120 14560
rect 4068 14408 4120 14414
rect 4068 14350 4120 14356
rect 4080 14006 4108 14350
rect 4068 14000 4120 14006
rect 4068 13942 4120 13948
rect 4160 13932 4212 13938
rect 4160 13874 4212 13880
rect 4172 13818 4200 13874
rect 4816 13870 4844 14962
rect 5000 14890 5028 15302
rect 5080 14952 5132 14958
rect 5080 14894 5132 14900
rect 4988 14884 5040 14890
rect 4988 14826 5040 14832
rect 5000 14414 5028 14826
rect 5092 14618 5120 14894
rect 5724 14816 5776 14822
rect 5724 14758 5776 14764
rect 5080 14612 5132 14618
rect 5080 14554 5132 14560
rect 4988 14408 5040 14414
rect 4988 14350 5040 14356
rect 5000 14278 5028 14350
rect 5264 14340 5316 14346
rect 5264 14282 5316 14288
rect 5356 14340 5408 14346
rect 5356 14282 5408 14288
rect 4988 14272 5040 14278
rect 4988 14214 5040 14220
rect 5276 14074 5304 14282
rect 5264 14068 5316 14074
rect 5264 14010 5316 14016
rect 5276 13938 5304 14010
rect 5264 13932 5316 13938
rect 5264 13874 5316 13880
rect 4080 13790 4200 13818
rect 4620 13864 4672 13870
rect 4620 13806 4672 13812
rect 4804 13864 4856 13870
rect 5368 13818 5396 14282
rect 5736 13938 5764 14758
rect 6092 14408 6144 14414
rect 6092 14350 6144 14356
rect 5816 14272 5868 14278
rect 5816 14214 5868 14220
rect 5828 13938 5856 14214
rect 6104 14006 6132 14350
rect 6472 14249 6500 18566
rect 6564 18426 6592 18702
rect 6552 18420 6604 18426
rect 6552 18362 6604 18368
rect 6564 17678 6592 18362
rect 6748 18222 6776 20703
rect 8214 20700 8522 20709
rect 8214 20698 8220 20700
rect 8276 20698 8300 20700
rect 8356 20698 8380 20700
rect 8436 20698 8460 20700
rect 8516 20698 8522 20700
rect 8276 20646 8278 20698
rect 8458 20646 8460 20698
rect 8214 20644 8220 20646
rect 8276 20644 8300 20646
rect 8356 20644 8380 20646
rect 8436 20644 8460 20646
rect 8516 20644 8522 20646
rect 8214 20635 8522 20644
rect 8760 20596 8812 20602
rect 8760 20538 8812 20544
rect 7380 20460 7432 20466
rect 7380 20402 7432 20408
rect 8576 20460 8628 20466
rect 8576 20402 8628 20408
rect 7012 19848 7064 19854
rect 7012 19790 7064 19796
rect 7024 19514 7052 19790
rect 7392 19786 7420 20402
rect 7472 20256 7524 20262
rect 7472 20198 7524 20204
rect 7380 19780 7432 19786
rect 7380 19722 7432 19728
rect 7012 19508 7064 19514
rect 7012 19450 7064 19456
rect 7484 19378 7512 20198
rect 8214 19612 8522 19621
rect 8214 19610 8220 19612
rect 8276 19610 8300 19612
rect 8356 19610 8380 19612
rect 8436 19610 8460 19612
rect 8516 19610 8522 19612
rect 8276 19558 8278 19610
rect 8458 19558 8460 19610
rect 8214 19556 8220 19558
rect 8276 19556 8300 19558
rect 8356 19556 8380 19558
rect 8436 19556 8460 19558
rect 8516 19556 8522 19558
rect 8214 19547 8522 19556
rect 8588 19378 8616 20402
rect 8772 19446 8800 20538
rect 9140 20466 9168 20946
rect 9416 20874 9444 21200
rect 9956 21004 10008 21010
rect 9956 20946 10008 20952
rect 9404 20868 9456 20874
rect 9404 20810 9456 20816
rect 9864 20528 9916 20534
rect 9864 20470 9916 20476
rect 9128 20460 9180 20466
rect 9128 20402 9180 20408
rect 9312 20460 9364 20466
rect 9312 20402 9364 20408
rect 9140 19938 9168 20402
rect 8956 19910 9168 19938
rect 8956 19854 8984 19910
rect 8944 19848 8996 19854
rect 8944 19790 8996 19796
rect 9128 19848 9180 19854
rect 9128 19790 9180 19796
rect 9324 19802 9352 20402
rect 9404 20256 9456 20262
rect 9404 20198 9456 20204
rect 9496 20256 9548 20262
rect 9496 20198 9548 20204
rect 9416 19990 9444 20198
rect 9404 19984 9456 19990
rect 9404 19926 9456 19932
rect 9508 19922 9536 20198
rect 9876 20058 9904 20470
rect 9864 20052 9916 20058
rect 9864 19994 9916 20000
rect 9496 19916 9548 19922
rect 9496 19858 9548 19864
rect 8760 19440 8812 19446
rect 8760 19382 8812 19388
rect 7104 19372 7156 19378
rect 7104 19314 7156 19320
rect 7472 19372 7524 19378
rect 7472 19314 7524 19320
rect 8576 19372 8628 19378
rect 8576 19314 8628 19320
rect 9036 19372 9088 19378
rect 9036 19314 9088 19320
rect 7116 18970 7144 19314
rect 7288 19168 7340 19174
rect 7288 19110 7340 19116
rect 7104 18964 7156 18970
rect 7104 18906 7156 18912
rect 6828 18896 6880 18902
rect 6828 18838 6880 18844
rect 6840 18290 6868 18838
rect 6920 18760 6972 18766
rect 6920 18702 6972 18708
rect 6828 18284 6880 18290
rect 6828 18226 6880 18232
rect 6736 18216 6788 18222
rect 6736 18158 6788 18164
rect 6552 17672 6604 17678
rect 6552 17614 6604 17620
rect 6932 15337 6960 18702
rect 7300 17746 7328 19110
rect 8588 18970 8616 19314
rect 9048 18970 9076 19314
rect 9140 19310 9168 19790
rect 9324 19774 9444 19802
rect 9416 19718 9444 19774
rect 9404 19712 9456 19718
rect 9404 19654 9456 19660
rect 9416 19514 9444 19654
rect 9404 19508 9456 19514
rect 9404 19450 9456 19456
rect 9968 19310 9996 20946
rect 11440 20806 11468 21200
rect 11428 20800 11480 20806
rect 11428 20742 11480 20748
rect 11980 20528 12032 20534
rect 11980 20470 12032 20476
rect 10048 20392 10100 20398
rect 10048 20334 10100 20340
rect 11152 20392 11204 20398
rect 11152 20334 11204 20340
rect 11244 20392 11296 20398
rect 11244 20334 11296 20340
rect 10060 19922 10088 20334
rect 10232 20324 10284 20330
rect 10232 20266 10284 20272
rect 10244 19922 10272 20266
rect 11164 19990 11192 20334
rect 11152 19984 11204 19990
rect 11152 19926 11204 19932
rect 10048 19916 10100 19922
rect 10048 19858 10100 19864
rect 10232 19916 10284 19922
rect 10232 19858 10284 19864
rect 10416 19916 10468 19922
rect 10416 19858 10468 19864
rect 10048 19440 10100 19446
rect 10048 19382 10100 19388
rect 9128 19304 9180 19310
rect 9128 19246 9180 19252
rect 9956 19304 10008 19310
rect 9956 19246 10008 19252
rect 9496 19236 9548 19242
rect 9496 19178 9548 19184
rect 8576 18964 8628 18970
rect 8576 18906 8628 18912
rect 9036 18964 9088 18970
rect 9036 18906 9088 18912
rect 7748 18828 7800 18834
rect 7748 18770 7800 18776
rect 7288 17740 7340 17746
rect 7288 17682 7340 17688
rect 7012 17672 7064 17678
rect 7012 17614 7064 17620
rect 7024 17270 7052 17614
rect 7012 17264 7064 17270
rect 7012 17206 7064 17212
rect 7024 16794 7052 17206
rect 7012 16788 7064 16794
rect 7012 16730 7064 16736
rect 7300 16590 7328 17682
rect 7564 17536 7616 17542
rect 7564 17478 7616 17484
rect 7576 17202 7604 17478
rect 7564 17196 7616 17202
rect 7564 17138 7616 17144
rect 7472 17128 7524 17134
rect 7472 17070 7524 17076
rect 7484 16658 7512 17070
rect 7472 16652 7524 16658
rect 7472 16594 7524 16600
rect 7288 16584 7340 16590
rect 7288 16526 7340 16532
rect 7380 16584 7432 16590
rect 7380 16526 7432 16532
rect 7656 16584 7708 16590
rect 7656 16526 7708 16532
rect 7392 16425 7420 16526
rect 7378 16416 7434 16425
rect 7378 16351 7434 16360
rect 7668 16250 7696 16526
rect 7760 16522 7788 18770
rect 7840 18692 7892 18698
rect 7840 18634 7892 18640
rect 7852 16998 7880 18634
rect 8214 18524 8522 18533
rect 8214 18522 8220 18524
rect 8276 18522 8300 18524
rect 8356 18522 8380 18524
rect 8436 18522 8460 18524
rect 8516 18522 8522 18524
rect 8276 18470 8278 18522
rect 8458 18470 8460 18522
rect 8214 18468 8220 18470
rect 8276 18468 8300 18470
rect 8356 18468 8380 18470
rect 8436 18468 8460 18470
rect 8516 18468 8522 18470
rect 8214 18459 8522 18468
rect 9404 17808 9456 17814
rect 9404 17750 9456 17756
rect 8576 17672 8628 17678
rect 8576 17614 8628 17620
rect 7932 17536 7984 17542
rect 7932 17478 7984 17484
rect 7944 17202 7972 17478
rect 8214 17436 8522 17445
rect 8214 17434 8220 17436
rect 8276 17434 8300 17436
rect 8356 17434 8380 17436
rect 8436 17434 8460 17436
rect 8516 17434 8522 17436
rect 8276 17382 8278 17434
rect 8458 17382 8460 17434
rect 8214 17380 8220 17382
rect 8276 17380 8300 17382
rect 8356 17380 8380 17382
rect 8436 17380 8460 17382
rect 8516 17380 8522 17382
rect 8214 17371 8522 17380
rect 7932 17196 7984 17202
rect 7932 17138 7984 17144
rect 8392 17196 8444 17202
rect 8392 17138 8444 17144
rect 7840 16992 7892 16998
rect 7840 16934 7892 16940
rect 7748 16516 7800 16522
rect 7748 16458 7800 16464
rect 7656 16244 7708 16250
rect 7656 16186 7708 16192
rect 7760 15978 7788 16458
rect 7748 15972 7800 15978
rect 7748 15914 7800 15920
rect 6918 15328 6974 15337
rect 6918 15263 6974 15272
rect 6828 15156 6880 15162
rect 6828 15098 6880 15104
rect 6840 14958 6868 15098
rect 6828 14952 6880 14958
rect 7104 14952 7156 14958
rect 6880 14912 6960 14940
rect 6828 14894 6880 14900
rect 6644 14408 6696 14414
rect 6644 14350 6696 14356
rect 6458 14240 6514 14249
rect 6458 14175 6514 14184
rect 6656 14074 6684 14350
rect 6828 14340 6880 14346
rect 6828 14282 6880 14288
rect 6644 14068 6696 14074
rect 6644 14010 6696 14016
rect 6840 14006 6868 14282
rect 6092 14000 6144 14006
rect 6092 13942 6144 13948
rect 6828 14000 6880 14006
rect 6828 13942 6880 13948
rect 5724 13932 5776 13938
rect 5724 13874 5776 13880
rect 5816 13932 5868 13938
rect 5816 13874 5868 13880
rect 4804 13806 4856 13812
rect 3976 13728 4028 13734
rect 3976 13670 4028 13676
rect 4080 13410 4108 13790
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4632 13462 4660 13806
rect 4620 13456 4672 13462
rect 3884 13388 3936 13394
rect 4080 13382 4200 13410
rect 4620 13398 4672 13404
rect 3884 13330 3936 13336
rect 3240 13320 3292 13326
rect 3240 13262 3292 13268
rect 3608 13320 3660 13326
rect 3608 13262 3660 13268
rect 3620 12850 3648 13262
rect 3608 12844 3660 12850
rect 3608 12786 3660 12792
rect 3896 12782 3924 13330
rect 4172 12850 4200 13382
rect 4160 12844 4212 12850
rect 4160 12786 4212 12792
rect 4632 12782 4660 13398
rect 4816 13394 4844 13806
rect 5276 13790 5396 13818
rect 4804 13388 4856 13394
rect 4804 13330 4856 13336
rect 5276 13326 5304 13790
rect 6460 13728 6512 13734
rect 6460 13670 6512 13676
rect 6472 13326 6500 13670
rect 4712 13320 4764 13326
rect 4712 13262 4764 13268
rect 5264 13320 5316 13326
rect 5264 13262 5316 13268
rect 5356 13320 5408 13326
rect 5356 13262 5408 13268
rect 5540 13320 5592 13326
rect 5540 13262 5592 13268
rect 6276 13320 6328 13326
rect 6276 13262 6328 13268
rect 6368 13320 6420 13326
rect 6368 13262 6420 13268
rect 6460 13320 6512 13326
rect 6460 13262 6512 13268
rect 4724 12850 4752 13262
rect 5276 12850 5304 13262
rect 5368 12918 5396 13262
rect 5356 12912 5408 12918
rect 5356 12854 5408 12860
rect 5552 12850 5580 13262
rect 6288 12850 6316 13262
rect 4712 12844 4764 12850
rect 4712 12786 4764 12792
rect 5264 12844 5316 12850
rect 5264 12786 5316 12792
rect 5540 12844 5592 12850
rect 5540 12786 5592 12792
rect 6276 12844 6328 12850
rect 6276 12786 6328 12792
rect 3884 12776 3936 12782
rect 3884 12718 3936 12724
rect 4620 12776 4672 12782
rect 4620 12718 4672 12724
rect 2412 12232 2464 12238
rect 2412 12174 2464 12180
rect 2688 12232 2740 12238
rect 2688 12174 2740 12180
rect 3424 12232 3476 12238
rect 3424 12174 3476 12180
rect 2424 11694 2452 12174
rect 2596 12096 2648 12102
rect 2596 12038 2648 12044
rect 2608 11830 2636 12038
rect 2596 11824 2648 11830
rect 2596 11766 2648 11772
rect 1492 11688 1544 11694
rect 1492 11630 1544 11636
rect 1952 11688 2004 11694
rect 1952 11630 2004 11636
rect 2412 11688 2464 11694
rect 2412 11630 2464 11636
rect 1306 10976 1362 10985
rect 1306 10911 1362 10920
rect 1320 10742 1348 10911
rect 1308 10736 1360 10742
rect 1308 10678 1360 10684
rect 1504 10062 1532 11630
rect 1964 11354 1992 11630
rect 1952 11348 2004 11354
rect 1952 11290 2004 11296
rect 2424 10674 2452 11630
rect 2700 10674 2728 12174
rect 3436 11558 3464 12174
rect 3424 11552 3476 11558
rect 3424 11494 3476 11500
rect 3332 11212 3384 11218
rect 3332 11154 3384 11160
rect 3240 11008 3292 11014
rect 3344 10996 3372 11154
rect 3436 11150 3464 11494
rect 3424 11144 3476 11150
rect 3424 11086 3476 11092
rect 3344 10968 3464 10996
rect 3240 10950 3292 10956
rect 3252 10810 3280 10950
rect 3240 10804 3292 10810
rect 3240 10746 3292 10752
rect 2412 10668 2464 10674
rect 2412 10610 2464 10616
rect 2688 10668 2740 10674
rect 2688 10610 2740 10616
rect 1492 10056 1544 10062
rect 1492 9998 1544 10004
rect 1306 8800 1362 8809
rect 1306 8735 1362 8744
rect 1320 8634 1348 8735
rect 1308 8628 1360 8634
rect 1308 8570 1360 8576
rect 1504 8430 1532 9998
rect 1768 9988 1820 9994
rect 1768 9930 1820 9936
rect 1780 9722 1808 9930
rect 1768 9716 1820 9722
rect 1768 9658 1820 9664
rect 2228 8968 2280 8974
rect 2228 8910 2280 8916
rect 1768 8832 1820 8838
rect 1768 8774 1820 8780
rect 1780 8566 1808 8774
rect 1768 8560 1820 8566
rect 1768 8502 1820 8508
rect 1492 8424 1544 8430
rect 1492 8366 1544 8372
rect 1504 6866 1532 8366
rect 2240 8090 2268 8910
rect 2228 8084 2280 8090
rect 2228 8026 2280 8032
rect 1860 7404 1912 7410
rect 1860 7346 1912 7352
rect 1492 6860 1544 6866
rect 1492 6802 1544 6808
rect 1504 5234 1532 6802
rect 1768 6724 1820 6730
rect 1768 6666 1820 6672
rect 1780 6458 1808 6666
rect 1768 6452 1820 6458
rect 1768 6394 1820 6400
rect 1492 5228 1544 5234
rect 1492 5170 1544 5176
rect 1504 4146 1532 5170
rect 1872 4622 1900 7346
rect 2424 6914 2452 10610
rect 2504 10464 2556 10470
rect 2504 10406 2556 10412
rect 2516 9994 2544 10406
rect 2504 9988 2556 9994
rect 2504 9930 2556 9936
rect 2504 7948 2556 7954
rect 2504 7890 2556 7896
rect 2516 7410 2544 7890
rect 2700 7886 2728 10610
rect 3240 10532 3292 10538
rect 3240 10474 3292 10480
rect 3252 9926 3280 10474
rect 3240 9920 3292 9926
rect 3240 9862 3292 9868
rect 3252 9722 3280 9862
rect 3240 9716 3292 9722
rect 3240 9658 3292 9664
rect 3436 9518 3464 10968
rect 3424 9512 3476 9518
rect 3424 9454 3476 9460
rect 3240 9036 3292 9042
rect 3240 8978 3292 8984
rect 2780 8560 2832 8566
rect 2780 8502 2832 8508
rect 2792 8022 2820 8502
rect 3252 8430 3280 8978
rect 3240 8424 3292 8430
rect 3240 8366 3292 8372
rect 2780 8016 2832 8022
rect 2780 7958 2832 7964
rect 3252 7886 3280 8366
rect 3436 7954 3464 9454
rect 3608 8968 3660 8974
rect 3608 8910 3660 8916
rect 3620 8634 3648 8910
rect 3896 8634 3924 12718
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 6380 12434 6408 13262
rect 6736 13252 6788 13258
rect 6736 13194 6788 13200
rect 6748 12918 6776 13194
rect 6736 12912 6788 12918
rect 6736 12854 6788 12860
rect 6104 12406 6408 12434
rect 4804 12300 4856 12306
rect 4804 12242 4856 12248
rect 3976 12096 4028 12102
rect 3976 12038 4028 12044
rect 3988 11762 4016 12038
rect 4540 11762 4752 11778
rect 3976 11756 4028 11762
rect 3976 11698 4028 11704
rect 4528 11756 4752 11762
rect 4580 11750 4752 11756
rect 4528 11698 4580 11704
rect 3988 11286 4016 11698
rect 4620 11620 4672 11626
rect 4620 11562 4672 11568
rect 4068 11552 4120 11558
rect 4068 11494 4120 11500
rect 3976 11280 4028 11286
rect 3976 11222 4028 11228
rect 3976 11144 4028 11150
rect 3976 11086 4028 11092
rect 3988 10674 4016 11086
rect 4080 11082 4108 11494
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4068 11076 4120 11082
rect 4068 11018 4120 11024
rect 4632 10674 4660 11562
rect 4724 11082 4752 11750
rect 4816 11354 4844 12242
rect 6000 12232 6052 12238
rect 6000 12174 6052 12180
rect 4896 12164 4948 12170
rect 4896 12106 4948 12112
rect 4804 11348 4856 11354
rect 4804 11290 4856 11296
rect 4712 11076 4764 11082
rect 4712 11018 4764 11024
rect 4724 10810 4752 11018
rect 4804 11008 4856 11014
rect 4804 10950 4856 10956
rect 4712 10804 4764 10810
rect 4712 10746 4764 10752
rect 3976 10668 4028 10674
rect 3976 10610 4028 10616
rect 4620 10668 4672 10674
rect 4620 10610 4672 10616
rect 3988 10198 4016 10610
rect 4068 10600 4120 10606
rect 4068 10542 4120 10548
rect 4080 10248 4108 10542
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4080 10220 4200 10248
rect 3976 10192 4028 10198
rect 3976 10134 4028 10140
rect 4172 9994 4200 10220
rect 4252 10124 4304 10130
rect 4252 10066 4304 10072
rect 4160 9988 4212 9994
rect 4160 9930 4212 9936
rect 4264 9654 4292 10066
rect 4436 9988 4488 9994
rect 4436 9930 4488 9936
rect 4448 9654 4476 9930
rect 4252 9648 4304 9654
rect 4252 9590 4304 9596
rect 4436 9648 4488 9654
rect 4436 9590 4488 9596
rect 4528 9580 4580 9586
rect 4528 9522 4580 9528
rect 4540 9466 4568 9522
rect 3976 9444 4028 9450
rect 4540 9438 4660 9466
rect 3976 9386 4028 9392
rect 3988 9110 4016 9386
rect 4068 9376 4120 9382
rect 4068 9318 4120 9324
rect 3976 9104 4028 9110
rect 3976 9046 4028 9052
rect 3608 8628 3660 8634
rect 3608 8570 3660 8576
rect 3884 8628 3936 8634
rect 3884 8570 3936 8576
rect 3620 8090 3648 8570
rect 4080 8498 4108 9318
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4632 9042 4660 9438
rect 4712 9444 4764 9450
rect 4712 9386 4764 9392
rect 4620 9036 4672 9042
rect 4620 8978 4672 8984
rect 4528 8832 4580 8838
rect 4528 8774 4580 8780
rect 4068 8492 4120 8498
rect 4068 8434 4120 8440
rect 4540 8362 4568 8774
rect 4528 8356 4580 8362
rect 4528 8298 4580 8304
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4632 8090 4660 8978
rect 4724 8974 4752 9386
rect 4712 8968 4764 8974
rect 4712 8910 4764 8916
rect 4712 8832 4764 8838
rect 4712 8774 4764 8780
rect 4724 8430 4752 8774
rect 4816 8498 4844 10950
rect 4908 10470 4936 12106
rect 5540 12096 5592 12102
rect 5540 12038 5592 12044
rect 5816 12096 5868 12102
rect 5816 12038 5868 12044
rect 5552 11218 5580 12038
rect 5828 11830 5856 12038
rect 5724 11824 5776 11830
rect 5724 11766 5776 11772
rect 5816 11824 5868 11830
rect 5816 11766 5868 11772
rect 5736 11286 5764 11766
rect 6012 11354 6040 12174
rect 6000 11348 6052 11354
rect 6000 11290 6052 11296
rect 5724 11280 5776 11286
rect 5724 11222 5776 11228
rect 5540 11212 5592 11218
rect 5540 11154 5592 11160
rect 4988 10804 5040 10810
rect 6104 10792 6132 12406
rect 6276 12164 6328 12170
rect 6276 12106 6328 12112
rect 6288 11354 6316 12106
rect 6932 11762 6960 14912
rect 7104 14894 7156 14900
rect 7116 14618 7144 14894
rect 7852 14822 7880 16934
rect 8404 16590 8432 17138
rect 8484 17128 8536 17134
rect 8484 17070 8536 17076
rect 8496 16674 8524 17070
rect 8588 16794 8616 17614
rect 9218 17368 9274 17377
rect 9218 17303 9274 17312
rect 9128 17196 9180 17202
rect 9128 17138 9180 17144
rect 9140 17066 9168 17138
rect 9128 17060 9180 17066
rect 9128 17002 9180 17008
rect 8576 16788 8628 16794
rect 8576 16730 8628 16736
rect 8496 16646 8800 16674
rect 8772 16590 8800 16646
rect 8392 16584 8444 16590
rect 8392 16526 8444 16532
rect 8760 16584 8812 16590
rect 8760 16526 8812 16532
rect 9140 16522 9168 17002
rect 8852 16516 8904 16522
rect 8852 16458 8904 16464
rect 9128 16516 9180 16522
rect 9128 16458 9180 16464
rect 8214 16348 8522 16357
rect 8214 16346 8220 16348
rect 8276 16346 8300 16348
rect 8356 16346 8380 16348
rect 8436 16346 8460 16348
rect 8516 16346 8522 16348
rect 8276 16294 8278 16346
rect 8458 16294 8460 16346
rect 8214 16292 8220 16294
rect 8276 16292 8300 16294
rect 8356 16292 8380 16294
rect 8436 16292 8460 16294
rect 8516 16292 8522 16294
rect 8214 16283 8522 16292
rect 8864 16250 8892 16458
rect 9232 16266 9260 17303
rect 9416 17202 9444 17750
rect 9404 17196 9456 17202
rect 9324 17156 9404 17184
rect 9324 16658 9352 17156
rect 9404 17138 9456 17144
rect 9508 17066 9536 19178
rect 9680 18964 9732 18970
rect 9680 18906 9732 18912
rect 9588 18828 9640 18834
rect 9588 18770 9640 18776
rect 9496 17060 9548 17066
rect 9496 17002 9548 17008
rect 9600 16658 9628 18770
rect 9692 18290 9720 18906
rect 10060 18902 10088 19382
rect 10428 19378 10456 19858
rect 10782 19816 10838 19825
rect 10782 19751 10838 19760
rect 10796 19446 10824 19751
rect 10876 19712 10928 19718
rect 10876 19654 10928 19660
rect 10784 19440 10836 19446
rect 10784 19382 10836 19388
rect 10888 19378 10916 19654
rect 11256 19514 11284 20334
rect 11992 20058 12020 20470
rect 12716 20392 12768 20398
rect 12716 20334 12768 20340
rect 12072 20324 12124 20330
rect 12072 20266 12124 20272
rect 12084 20058 12112 20266
rect 12728 20262 12756 20334
rect 12716 20256 12768 20262
rect 12716 20198 12768 20204
rect 12214 20156 12522 20165
rect 12214 20154 12220 20156
rect 12276 20154 12300 20156
rect 12356 20154 12380 20156
rect 12436 20154 12460 20156
rect 12516 20154 12522 20156
rect 12276 20102 12278 20154
rect 12458 20102 12460 20154
rect 12214 20100 12220 20102
rect 12276 20100 12300 20102
rect 12356 20100 12380 20102
rect 12436 20100 12460 20102
rect 12516 20100 12522 20102
rect 12214 20091 12522 20100
rect 11980 20052 12032 20058
rect 11980 19994 12032 20000
rect 12072 20052 12124 20058
rect 12072 19994 12124 20000
rect 11992 19854 12020 19994
rect 11612 19848 11664 19854
rect 11612 19790 11664 19796
rect 11980 19848 12032 19854
rect 11980 19790 12032 19796
rect 11428 19780 11480 19786
rect 11428 19722 11480 19728
rect 11244 19508 11296 19514
rect 11244 19450 11296 19456
rect 10416 19372 10468 19378
rect 10416 19314 10468 19320
rect 10876 19372 10928 19378
rect 10876 19314 10928 19320
rect 11060 19372 11112 19378
rect 11060 19314 11112 19320
rect 10888 19242 10916 19314
rect 10876 19236 10928 19242
rect 10876 19178 10928 19184
rect 10888 18970 10916 19178
rect 10508 18964 10560 18970
rect 10508 18906 10560 18912
rect 10876 18964 10928 18970
rect 10876 18906 10928 18912
rect 10048 18896 10100 18902
rect 10048 18838 10100 18844
rect 10140 18760 10192 18766
rect 10140 18702 10192 18708
rect 9680 18284 9732 18290
rect 9680 18226 9732 18232
rect 10152 18222 10180 18702
rect 10520 18358 10548 18906
rect 10876 18420 10928 18426
rect 10876 18362 10928 18368
rect 10508 18352 10560 18358
rect 10336 18312 10508 18340
rect 10140 18216 10192 18222
rect 10140 18158 10192 18164
rect 9864 18148 9916 18154
rect 9864 18090 9916 18096
rect 9772 17672 9824 17678
rect 9772 17614 9824 17620
rect 9680 17196 9732 17202
rect 9680 17138 9732 17144
rect 9312 16652 9364 16658
rect 9312 16594 9364 16600
rect 9588 16652 9640 16658
rect 9588 16594 9640 16600
rect 9496 16448 9548 16454
rect 9496 16390 9548 16396
rect 8852 16244 8904 16250
rect 8852 16186 8904 16192
rect 9140 16238 9260 16266
rect 9508 16250 9536 16390
rect 9496 16244 9548 16250
rect 9140 16114 9168 16238
rect 9496 16186 9548 16192
rect 8300 16108 8352 16114
rect 8300 16050 8352 16056
rect 9128 16108 9180 16114
rect 9128 16050 9180 16056
rect 9220 16108 9272 16114
rect 9220 16050 9272 16056
rect 9312 16108 9364 16114
rect 9312 16050 9364 16056
rect 8024 15904 8076 15910
rect 8024 15846 8076 15852
rect 8036 15502 8064 15846
rect 8024 15496 8076 15502
rect 8024 15438 8076 15444
rect 8312 15434 8340 16050
rect 8668 15564 8720 15570
rect 8668 15506 8720 15512
rect 8576 15496 8628 15502
rect 8576 15438 8628 15444
rect 8300 15428 8352 15434
rect 8300 15370 8352 15376
rect 8116 15360 8168 15366
rect 8116 15302 8168 15308
rect 8128 15094 8156 15302
rect 8214 15260 8522 15269
rect 8214 15258 8220 15260
rect 8276 15258 8300 15260
rect 8356 15258 8380 15260
rect 8436 15258 8460 15260
rect 8516 15258 8522 15260
rect 8276 15206 8278 15258
rect 8458 15206 8460 15258
rect 8214 15204 8220 15206
rect 8276 15204 8300 15206
rect 8356 15204 8380 15206
rect 8436 15204 8460 15206
rect 8516 15204 8522 15206
rect 8214 15195 8522 15204
rect 8588 15162 8616 15438
rect 8576 15156 8628 15162
rect 8576 15098 8628 15104
rect 8116 15088 8168 15094
rect 8116 15030 8168 15036
rect 7840 14816 7892 14822
rect 7840 14758 7892 14764
rect 8680 14618 8708 15506
rect 8852 15428 8904 15434
rect 8852 15370 8904 15376
rect 7104 14612 7156 14618
rect 7104 14554 7156 14560
rect 8668 14612 8720 14618
rect 8668 14554 8720 14560
rect 8576 14476 8628 14482
rect 8576 14418 8628 14424
rect 7288 14408 7340 14414
rect 7288 14350 7340 14356
rect 7104 13796 7156 13802
rect 7104 13738 7156 13744
rect 7116 13326 7144 13738
rect 7300 13394 7328 14350
rect 7748 14272 7800 14278
rect 7748 14214 7800 14220
rect 7760 14074 7788 14214
rect 8214 14172 8522 14181
rect 8214 14170 8220 14172
rect 8276 14170 8300 14172
rect 8356 14170 8380 14172
rect 8436 14170 8460 14172
rect 8516 14170 8522 14172
rect 8276 14118 8278 14170
rect 8458 14118 8460 14170
rect 8214 14116 8220 14118
rect 8276 14116 8300 14118
rect 8356 14116 8380 14118
rect 8436 14116 8460 14118
rect 8516 14116 8522 14118
rect 8214 14107 8522 14116
rect 7748 14068 7800 14074
rect 7748 14010 7800 14016
rect 8300 14000 8352 14006
rect 8352 13948 8524 13954
rect 8300 13942 8524 13948
rect 8312 13938 8524 13942
rect 8588 13938 8616 14418
rect 8864 14414 8892 15370
rect 9140 15026 9168 16050
rect 9232 15706 9260 16050
rect 9220 15700 9272 15706
rect 9220 15642 9272 15648
rect 9128 15020 9180 15026
rect 9128 14962 9180 14968
rect 9232 14414 9260 15642
rect 9324 14890 9352 16050
rect 9600 15978 9628 16594
rect 9692 16522 9720 17138
rect 9680 16516 9732 16522
rect 9680 16458 9732 16464
rect 9784 16425 9812 17614
rect 9876 17202 9904 18090
rect 10152 17610 10180 18158
rect 10336 17882 10364 18312
rect 10508 18294 10560 18300
rect 10414 18184 10470 18193
rect 10414 18119 10470 18128
rect 10324 17876 10376 17882
rect 10324 17818 10376 17824
rect 10232 17740 10284 17746
rect 10232 17682 10284 17688
rect 10140 17604 10192 17610
rect 10140 17546 10192 17552
rect 10152 17513 10180 17546
rect 10138 17504 10194 17513
rect 10138 17439 10194 17448
rect 10244 17241 10272 17682
rect 10230 17232 10286 17241
rect 9864 17196 9916 17202
rect 9864 17138 9916 17144
rect 9956 17196 10008 17202
rect 10140 17196 10192 17202
rect 9956 17138 10008 17144
rect 10060 17156 10140 17184
rect 9876 17105 9904 17138
rect 9862 17096 9918 17105
rect 9968 17066 9996 17138
rect 9862 17031 9918 17040
rect 9956 17060 10008 17066
rect 9956 17002 10008 17008
rect 10060 16998 10088 17156
rect 10230 17167 10286 17176
rect 10140 17138 10192 17144
rect 10232 17060 10284 17066
rect 10232 17002 10284 17008
rect 10048 16992 10100 16998
rect 10048 16934 10100 16940
rect 10140 16584 10192 16590
rect 10140 16526 10192 16532
rect 9770 16416 9826 16425
rect 9770 16351 9826 16360
rect 9588 15972 9640 15978
rect 9588 15914 9640 15920
rect 10048 15972 10100 15978
rect 10048 15914 10100 15920
rect 9404 15496 9456 15502
rect 9404 15438 9456 15444
rect 9312 14884 9364 14890
rect 9312 14826 9364 14832
rect 9324 14482 9352 14826
rect 9312 14476 9364 14482
rect 9312 14418 9364 14424
rect 8852 14408 8904 14414
rect 8852 14350 8904 14356
rect 9220 14408 9272 14414
rect 9220 14350 9272 14356
rect 7472 13932 7524 13938
rect 8312 13932 8536 13938
rect 8312 13926 8484 13932
rect 7472 13874 7524 13880
rect 8484 13874 8536 13880
rect 8576 13932 8628 13938
rect 8576 13874 8628 13880
rect 7484 13530 7512 13874
rect 7564 13864 7616 13870
rect 7564 13806 7616 13812
rect 7472 13524 7524 13530
rect 7472 13466 7524 13472
rect 7288 13388 7340 13394
rect 7288 13330 7340 13336
rect 7104 13320 7156 13326
rect 7104 13262 7156 13268
rect 7576 13258 7604 13806
rect 8496 13802 8524 13874
rect 8484 13796 8536 13802
rect 8484 13738 8536 13744
rect 8496 13326 8524 13738
rect 8588 13530 8616 13874
rect 8760 13728 8812 13734
rect 8760 13670 8812 13676
rect 8576 13524 8628 13530
rect 8576 13466 8628 13472
rect 8772 13394 8800 13670
rect 8760 13388 8812 13394
rect 8760 13330 8812 13336
rect 8484 13320 8536 13326
rect 8484 13262 8536 13268
rect 7012 13252 7064 13258
rect 7012 13194 7064 13200
rect 7564 13252 7616 13258
rect 7564 13194 7616 13200
rect 7024 12782 7052 13194
rect 8214 13084 8522 13093
rect 8214 13082 8220 13084
rect 8276 13082 8300 13084
rect 8356 13082 8380 13084
rect 8436 13082 8460 13084
rect 8516 13082 8522 13084
rect 8276 13030 8278 13082
rect 8458 13030 8460 13082
rect 8214 13028 8220 13030
rect 8276 13028 8300 13030
rect 8356 13028 8380 13030
rect 8436 13028 8460 13030
rect 8516 13028 8522 13030
rect 8214 13019 8522 13028
rect 8864 12986 8892 14350
rect 8944 14340 8996 14346
rect 8944 14282 8996 14288
rect 9036 14340 9088 14346
rect 9036 14282 9088 14288
rect 8956 13938 8984 14282
rect 8944 13932 8996 13938
rect 8944 13874 8996 13880
rect 9048 13802 9076 14282
rect 9128 14272 9180 14278
rect 9128 14214 9180 14220
rect 9140 14006 9168 14214
rect 9128 14000 9180 14006
rect 9128 13942 9180 13948
rect 9036 13796 9088 13802
rect 9036 13738 9088 13744
rect 9220 13320 9272 13326
rect 9220 13262 9272 13268
rect 9232 12986 9260 13262
rect 8852 12980 8904 12986
rect 8852 12922 8904 12928
rect 9220 12980 9272 12986
rect 9220 12922 9272 12928
rect 9416 12918 9444 15438
rect 9600 15434 9628 15914
rect 9864 15904 9916 15910
rect 9916 15852 9996 15858
rect 9864 15846 9996 15852
rect 9876 15830 9996 15846
rect 9772 15632 9824 15638
rect 9772 15574 9824 15580
rect 9588 15428 9640 15434
rect 9588 15370 9640 15376
rect 9496 13932 9548 13938
rect 9496 13874 9548 13880
rect 9404 12912 9456 12918
rect 9404 12854 9456 12860
rect 7012 12776 7064 12782
rect 7012 12718 7064 12724
rect 9508 12714 9536 13874
rect 9600 13326 9628 15370
rect 9680 14952 9732 14958
rect 9680 14894 9732 14900
rect 9692 14618 9720 14894
rect 9680 14612 9732 14618
rect 9680 14554 9732 14560
rect 9692 13326 9720 14554
rect 9784 14482 9812 15574
rect 9864 15088 9916 15094
rect 9864 15030 9916 15036
rect 9876 14618 9904 15030
rect 9864 14612 9916 14618
rect 9864 14554 9916 14560
rect 9772 14476 9824 14482
rect 9772 14418 9824 14424
rect 9876 14006 9904 14554
rect 9864 14000 9916 14006
rect 9864 13942 9916 13948
rect 9968 13852 9996 15830
rect 10060 15162 10088 15914
rect 10152 15366 10180 16526
rect 10244 16046 10272 17002
rect 10232 16040 10284 16046
rect 10232 15982 10284 15988
rect 10336 15910 10364 17818
rect 10428 17678 10456 18119
rect 10692 18080 10744 18086
rect 10692 18022 10744 18028
rect 10600 17808 10652 17814
rect 10600 17750 10652 17756
rect 10612 17678 10640 17750
rect 10416 17672 10468 17678
rect 10600 17672 10652 17678
rect 10416 17614 10468 17620
rect 10520 17632 10600 17660
rect 10428 16697 10456 17614
rect 10520 17202 10548 17632
rect 10704 17649 10732 18022
rect 10888 17785 10916 18362
rect 10966 18320 11022 18329
rect 10966 18255 11022 18264
rect 10874 17776 10930 17785
rect 10874 17711 10930 17720
rect 10980 17678 11008 18255
rect 10968 17672 11020 17678
rect 10600 17614 10652 17620
rect 10690 17640 10746 17649
rect 10968 17614 11020 17620
rect 10690 17575 10746 17584
rect 10784 17604 10836 17610
rect 10598 17232 10654 17241
rect 10508 17196 10560 17202
rect 10598 17167 10600 17176
rect 10508 17138 10560 17144
rect 10652 17167 10654 17176
rect 10600 17138 10652 17144
rect 10414 16688 10470 16697
rect 10414 16623 10470 16632
rect 10324 15904 10376 15910
rect 10324 15846 10376 15852
rect 10428 15638 10456 16623
rect 10508 16584 10560 16590
rect 10508 16526 10560 16532
rect 10520 16182 10548 16526
rect 10508 16176 10560 16182
rect 10508 16118 10560 16124
rect 10704 16114 10732 17575
rect 10784 17546 10836 17552
rect 10796 16250 10824 17546
rect 10876 17536 10928 17542
rect 10876 17478 10928 17484
rect 10888 17338 10916 17478
rect 10876 17332 10928 17338
rect 10876 17274 10928 17280
rect 10980 17218 11008 17614
rect 10888 17190 11008 17218
rect 10888 16590 10916 17190
rect 10968 17060 11020 17066
rect 10968 17002 11020 17008
rect 10876 16584 10928 16590
rect 10876 16526 10928 16532
rect 10784 16244 10836 16250
rect 10784 16186 10836 16192
rect 10692 16108 10744 16114
rect 10692 16050 10744 16056
rect 10416 15632 10468 15638
rect 10416 15574 10468 15580
rect 10232 15564 10284 15570
rect 10232 15506 10284 15512
rect 10140 15360 10192 15366
rect 10140 15302 10192 15308
rect 10048 15156 10100 15162
rect 10048 15098 10100 15104
rect 10244 15026 10272 15506
rect 10324 15428 10376 15434
rect 10324 15370 10376 15376
rect 10048 15020 10100 15026
rect 10048 14962 10100 14968
rect 10232 15020 10284 15026
rect 10232 14962 10284 14968
rect 9876 13824 9996 13852
rect 9876 13326 9904 13824
rect 9588 13320 9640 13326
rect 9588 13262 9640 13268
rect 9680 13320 9732 13326
rect 9680 13262 9732 13268
rect 9864 13320 9916 13326
rect 9864 13262 9916 13268
rect 9692 13002 9720 13262
rect 9600 12974 9720 13002
rect 9496 12708 9548 12714
rect 9496 12650 9548 12656
rect 8576 12640 8628 12646
rect 8576 12582 8628 12588
rect 7012 12368 7064 12374
rect 7012 12310 7064 12316
rect 6920 11756 6972 11762
rect 6920 11698 6972 11704
rect 6828 11688 6880 11694
rect 6828 11630 6880 11636
rect 6736 11620 6788 11626
rect 6736 11562 6788 11568
rect 6276 11348 6328 11354
rect 6276 11290 6328 11296
rect 6552 11144 6604 11150
rect 6552 11086 6604 11092
rect 4988 10746 5040 10752
rect 6012 10764 6132 10792
rect 4896 10464 4948 10470
rect 4896 10406 4948 10412
rect 5000 9450 5028 10746
rect 5816 10668 5868 10674
rect 5816 10610 5868 10616
rect 5540 10600 5592 10606
rect 5540 10542 5592 10548
rect 5448 10464 5500 10470
rect 5448 10406 5500 10412
rect 5460 10062 5488 10406
rect 5448 10056 5500 10062
rect 5448 9998 5500 10004
rect 5552 9994 5580 10542
rect 5632 10464 5684 10470
rect 5632 10406 5684 10412
rect 5724 10464 5776 10470
rect 5724 10406 5776 10412
rect 5540 9988 5592 9994
rect 5540 9930 5592 9936
rect 5356 9920 5408 9926
rect 5356 9862 5408 9868
rect 5368 9586 5396 9862
rect 5356 9580 5408 9586
rect 5356 9522 5408 9528
rect 5552 9466 5580 9930
rect 5644 9586 5672 10406
rect 5736 10198 5764 10406
rect 5724 10192 5776 10198
rect 5724 10134 5776 10140
rect 5828 10062 5856 10610
rect 5816 10056 5868 10062
rect 5816 9998 5868 10004
rect 5908 10056 5960 10062
rect 5908 9998 5960 10004
rect 5828 9602 5856 9998
rect 5920 9722 5948 9998
rect 5908 9716 5960 9722
rect 5908 9658 5960 9664
rect 5828 9586 5948 9602
rect 5632 9580 5684 9586
rect 5632 9522 5684 9528
rect 5724 9580 5776 9586
rect 5828 9580 5960 9586
rect 5828 9574 5908 9580
rect 5724 9522 5776 9528
rect 5908 9522 5960 9528
rect 5736 9466 5764 9522
rect 4988 9444 5040 9450
rect 5552 9438 5764 9466
rect 4988 9386 5040 9392
rect 4988 8968 5040 8974
rect 6012 8922 6040 10764
rect 6092 10668 6144 10674
rect 6092 10610 6144 10616
rect 6104 10130 6132 10610
rect 6184 10600 6236 10606
rect 6184 10542 6236 10548
rect 6460 10600 6512 10606
rect 6460 10542 6512 10548
rect 6092 10124 6144 10130
rect 6092 10066 6144 10072
rect 6196 10062 6224 10542
rect 6368 10464 6420 10470
rect 6368 10406 6420 10412
rect 6184 10056 6236 10062
rect 6184 9998 6236 10004
rect 6276 10056 6328 10062
rect 6276 9998 6328 10004
rect 6092 9988 6144 9994
rect 6092 9930 6144 9936
rect 6104 9654 6132 9930
rect 6196 9897 6224 9998
rect 6182 9888 6238 9897
rect 6182 9823 6238 9832
rect 6092 9648 6144 9654
rect 6092 9590 6144 9596
rect 6288 9586 6316 9998
rect 6276 9580 6328 9586
rect 6276 9522 6328 9528
rect 4988 8910 5040 8916
rect 4896 8832 4948 8838
rect 4896 8774 4948 8780
rect 4804 8492 4856 8498
rect 4804 8434 4856 8440
rect 4908 8430 4936 8774
rect 4712 8424 4764 8430
rect 4712 8366 4764 8372
rect 4896 8424 4948 8430
rect 4896 8366 4948 8372
rect 3608 8084 3660 8090
rect 3608 8026 3660 8032
rect 4620 8084 4672 8090
rect 4620 8026 4672 8032
rect 3424 7948 3476 7954
rect 3424 7890 3476 7896
rect 2688 7880 2740 7886
rect 2688 7822 2740 7828
rect 3240 7880 3292 7886
rect 3240 7822 3292 7828
rect 2700 7410 2728 7822
rect 2504 7404 2556 7410
rect 2504 7346 2556 7352
rect 2688 7404 2740 7410
rect 2688 7346 2740 7352
rect 2780 7200 2832 7206
rect 2780 7142 2832 7148
rect 2424 6886 2544 6914
rect 2516 5710 2544 6886
rect 2792 6730 2820 7142
rect 2780 6724 2832 6730
rect 2780 6666 2832 6672
rect 3148 6656 3200 6662
rect 3148 6598 3200 6604
rect 3330 6624 3386 6633
rect 3160 6458 3188 6598
rect 3330 6559 3386 6568
rect 3148 6452 3200 6458
rect 3148 6394 3200 6400
rect 2872 6112 2924 6118
rect 2872 6054 2924 6060
rect 2780 5840 2832 5846
rect 2780 5782 2832 5788
rect 2504 5704 2556 5710
rect 2504 5646 2556 5652
rect 2044 5568 2096 5574
rect 2044 5510 2096 5516
rect 2056 5302 2084 5510
rect 2044 5296 2096 5302
rect 2044 5238 2096 5244
rect 2516 4690 2544 5646
rect 2792 5302 2820 5782
rect 2884 5710 2912 6054
rect 3344 5710 3372 6559
rect 3436 6254 3464 7890
rect 4068 7880 4120 7886
rect 4068 7822 4120 7828
rect 4080 7410 4108 7822
rect 4436 7744 4488 7750
rect 4436 7686 4488 7692
rect 4448 7546 4476 7686
rect 4436 7540 4488 7546
rect 4436 7482 4488 7488
rect 4068 7404 4120 7410
rect 4068 7346 4120 7352
rect 4080 7002 4108 7346
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4068 6996 4120 7002
rect 4068 6938 4120 6944
rect 3424 6248 3476 6254
rect 3424 6190 3476 6196
rect 3976 6248 4028 6254
rect 3976 6190 4028 6196
rect 2872 5704 2924 5710
rect 2872 5646 2924 5652
rect 3332 5704 3384 5710
rect 3332 5646 3384 5652
rect 3516 5704 3568 5710
rect 3516 5646 3568 5652
rect 2780 5296 2832 5302
rect 2780 5238 2832 5244
rect 2504 4684 2556 4690
rect 2504 4626 2556 4632
rect 1860 4616 1912 4622
rect 1860 4558 1912 4564
rect 1492 4140 1544 4146
rect 1492 4082 1544 4088
rect 1504 2854 1532 4082
rect 1952 4072 2004 4078
rect 1952 4014 2004 4020
rect 1964 3738 1992 4014
rect 1952 3732 2004 3738
rect 1952 3674 2004 3680
rect 2516 3466 2544 4626
rect 2884 3534 2912 5646
rect 3240 5636 3292 5642
rect 3240 5578 3292 5584
rect 3148 5568 3200 5574
rect 3054 5536 3110 5545
rect 3148 5510 3200 5516
rect 3054 5471 3110 5480
rect 3068 4690 3096 5471
rect 3056 4684 3108 4690
rect 3056 4626 3108 4632
rect 2964 4208 3016 4214
rect 2964 4150 3016 4156
rect 2976 3738 3004 4150
rect 3068 4010 3096 4626
rect 3160 4622 3188 5510
rect 3252 5370 3280 5578
rect 3240 5364 3292 5370
rect 3240 5306 3292 5312
rect 3344 5234 3372 5646
rect 3528 5352 3556 5646
rect 3608 5364 3660 5370
rect 3528 5324 3608 5352
rect 3332 5228 3384 5234
rect 3332 5170 3384 5176
rect 3528 5166 3556 5324
rect 3608 5306 3660 5312
rect 3792 5296 3844 5302
rect 3792 5238 3844 5244
rect 3516 5160 3568 5166
rect 3516 5102 3568 5108
rect 3528 4690 3556 5102
rect 3804 4826 3832 5238
rect 3988 5166 4016 6190
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4724 5846 4752 8366
rect 4908 7886 4936 8366
rect 4896 7880 4948 7886
rect 4896 7822 4948 7828
rect 4896 7744 4948 7750
rect 5000 7721 5028 8910
rect 5920 8894 6040 8922
rect 5080 8560 5132 8566
rect 5080 8502 5132 8508
rect 4896 7686 4948 7692
rect 4986 7712 5042 7721
rect 4908 7478 4936 7686
rect 4986 7647 5042 7656
rect 4896 7472 4948 7478
rect 4896 7414 4948 7420
rect 4804 6724 4856 6730
rect 4804 6666 4856 6672
rect 4816 6390 4844 6666
rect 4896 6656 4948 6662
rect 4896 6598 4948 6604
rect 4908 6390 4936 6598
rect 4804 6384 4856 6390
rect 4804 6326 4856 6332
rect 4896 6384 4948 6390
rect 4896 6326 4948 6332
rect 4712 5840 4764 5846
rect 4712 5782 4764 5788
rect 4712 5704 4764 5710
rect 4764 5664 4844 5692
rect 4712 5646 4764 5652
rect 4816 5302 4844 5664
rect 4804 5296 4856 5302
rect 4804 5238 4856 5244
rect 4528 5228 4580 5234
rect 4528 5170 4580 5176
rect 4712 5228 4764 5234
rect 4712 5170 4764 5176
rect 4896 5228 4948 5234
rect 4896 5170 4948 5176
rect 4988 5228 5040 5234
rect 4988 5170 5040 5176
rect 3976 5160 4028 5166
rect 3976 5102 4028 5108
rect 4540 5114 4568 5170
rect 3792 4820 3844 4826
rect 3792 4762 3844 4768
rect 3516 4684 3568 4690
rect 3516 4626 3568 4632
rect 3148 4616 3200 4622
rect 3148 4558 3200 4564
rect 3700 4480 3752 4486
rect 3700 4422 3752 4428
rect 3712 4146 3740 4422
rect 3700 4140 3752 4146
rect 3700 4082 3752 4088
rect 3056 4004 3108 4010
rect 3056 3946 3108 3952
rect 2964 3732 3016 3738
rect 2964 3674 3016 3680
rect 2872 3528 2924 3534
rect 2872 3470 2924 3476
rect 2504 3460 2556 3466
rect 2504 3402 2556 3408
rect 2516 3058 2544 3402
rect 2884 3398 2912 3470
rect 2872 3392 2924 3398
rect 2872 3334 2924 3340
rect 3608 3392 3660 3398
rect 3608 3334 3660 3340
rect 3620 3058 3648 3334
rect 2504 3052 2556 3058
rect 2504 2994 2556 3000
rect 3608 3052 3660 3058
rect 3608 2994 3660 3000
rect 3988 2854 4016 5102
rect 4540 5086 4660 5114
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4160 4684 4212 4690
rect 4160 4626 4212 4632
rect 4172 4282 4200 4626
rect 4632 4282 4660 5086
rect 4160 4276 4212 4282
rect 4160 4218 4212 4224
rect 4620 4276 4672 4282
rect 4620 4218 4672 4224
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4620 3392 4672 3398
rect 4620 3334 4672 3340
rect 4068 2916 4120 2922
rect 4068 2858 4120 2864
rect 1492 2848 1544 2854
rect 1492 2790 1544 2796
rect 2872 2848 2924 2854
rect 2872 2790 2924 2796
rect 3976 2848 4028 2854
rect 3976 2790 4028 2796
rect 202 2544 258 2553
rect 2884 2514 2912 2790
rect 4080 2530 4108 2858
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 202 2479 258 2488
rect 2872 2508 2924 2514
rect 4080 2502 4200 2530
rect 2872 2450 2924 2456
rect 2884 1970 2912 2450
rect 3148 2304 3200 2310
rect 3148 2246 3200 2252
rect 3160 2038 3188 2246
rect 4172 2038 4200 2502
rect 4632 2378 4660 3334
rect 4724 3194 4752 5170
rect 4908 4826 4936 5170
rect 4896 4820 4948 4826
rect 4896 4762 4948 4768
rect 4804 4616 4856 4622
rect 4804 4558 4856 4564
rect 4816 4146 4844 4558
rect 5000 4146 5028 5170
rect 5092 5098 5120 8502
rect 5172 8492 5224 8498
rect 5172 8434 5224 8440
rect 5184 8022 5212 8434
rect 5540 8356 5592 8362
rect 5540 8298 5592 8304
rect 5172 8016 5224 8022
rect 5172 7958 5224 7964
rect 5184 7410 5212 7958
rect 5552 7818 5580 8298
rect 5816 7880 5868 7886
rect 5816 7822 5868 7828
rect 5540 7812 5592 7818
rect 5540 7754 5592 7760
rect 5172 7404 5224 7410
rect 5552 7392 5580 7754
rect 5724 7744 5776 7750
rect 5724 7686 5776 7692
rect 5736 7546 5764 7686
rect 5828 7546 5856 7822
rect 5724 7540 5776 7546
rect 5724 7482 5776 7488
rect 5816 7540 5868 7546
rect 5816 7482 5868 7488
rect 5552 7364 5672 7392
rect 5172 7346 5224 7352
rect 5540 7268 5592 7274
rect 5540 7210 5592 7216
rect 5552 6866 5580 7210
rect 5172 6860 5224 6866
rect 5172 6802 5224 6808
rect 5540 6860 5592 6866
rect 5540 6802 5592 6808
rect 5184 6322 5212 6802
rect 5644 6798 5672 7364
rect 5632 6792 5684 6798
rect 5632 6734 5684 6740
rect 5736 6730 5764 7482
rect 5724 6724 5776 6730
rect 5724 6666 5776 6672
rect 5448 6656 5500 6662
rect 5448 6598 5500 6604
rect 5460 6322 5488 6598
rect 5172 6316 5224 6322
rect 5172 6258 5224 6264
rect 5448 6316 5500 6322
rect 5448 6258 5500 6264
rect 5184 5914 5212 6258
rect 5540 6248 5592 6254
rect 5540 6190 5592 6196
rect 5172 5908 5224 5914
rect 5172 5850 5224 5856
rect 5172 5704 5224 5710
rect 5172 5646 5224 5652
rect 5264 5704 5316 5710
rect 5264 5646 5316 5652
rect 5080 5092 5132 5098
rect 5080 5034 5132 5040
rect 5078 4448 5134 4457
rect 5078 4383 5134 4392
rect 4804 4140 4856 4146
rect 4804 4082 4856 4088
rect 4988 4140 5040 4146
rect 4988 4082 5040 4088
rect 4804 3936 4856 3942
rect 4804 3878 4856 3884
rect 4816 3602 4844 3878
rect 4804 3596 4856 3602
rect 4804 3538 4856 3544
rect 4712 3188 4764 3194
rect 4712 3130 4764 3136
rect 4804 2984 4856 2990
rect 4804 2926 4856 2932
rect 4988 2984 5040 2990
rect 4988 2926 5040 2932
rect 4816 2774 4844 2926
rect 4816 2746 4936 2774
rect 4436 2372 4488 2378
rect 4436 2314 4488 2320
rect 4620 2372 4672 2378
rect 4620 2314 4672 2320
rect 4448 2038 4476 2314
rect 4908 2106 4936 2746
rect 4896 2100 4948 2106
rect 4896 2042 4948 2048
rect 3148 2032 3200 2038
rect 3148 1974 3200 1980
rect 4160 2032 4212 2038
rect 4160 1974 4212 1980
rect 4436 2032 4488 2038
rect 4436 1974 4488 1980
rect 2872 1964 2924 1970
rect 2872 1906 2924 1912
rect 848 1420 900 1426
rect 848 1362 900 1368
rect 860 1329 888 1362
rect 2884 1358 2912 1906
rect 4896 1896 4948 1902
rect 4896 1838 4948 1844
rect 4214 1660 4522 1669
rect 4214 1658 4220 1660
rect 4276 1658 4300 1660
rect 4356 1658 4380 1660
rect 4436 1658 4460 1660
rect 4516 1658 4522 1660
rect 4276 1606 4278 1658
rect 4458 1606 4460 1658
rect 4214 1604 4220 1606
rect 4276 1604 4300 1606
rect 4356 1604 4380 1606
rect 4436 1604 4460 1606
rect 4516 1604 4522 1606
rect 4214 1595 4522 1604
rect 4908 1358 4936 1838
rect 5000 1562 5028 2926
rect 5092 1834 5120 4383
rect 5184 3194 5212 5646
rect 5276 4758 5304 5646
rect 5552 4758 5580 6190
rect 5920 5574 5948 8894
rect 6000 8832 6052 8838
rect 6000 8774 6052 8780
rect 6012 8430 6040 8774
rect 6000 8424 6052 8430
rect 6000 8366 6052 8372
rect 6380 8090 6408 10406
rect 6472 10266 6500 10542
rect 6564 10538 6592 11086
rect 6644 10736 6696 10742
rect 6644 10678 6696 10684
rect 6552 10532 6604 10538
rect 6552 10474 6604 10480
rect 6460 10260 6512 10266
rect 6460 10202 6512 10208
rect 6472 10130 6500 10202
rect 6460 10124 6512 10130
rect 6460 10066 6512 10072
rect 6656 9926 6684 10678
rect 6552 9920 6604 9926
rect 6552 9862 6604 9868
rect 6644 9920 6696 9926
rect 6644 9862 6696 9868
rect 6564 9654 6592 9862
rect 6748 9738 6776 11562
rect 6840 11150 6868 11630
rect 7024 11150 7052 12310
rect 8214 11996 8522 12005
rect 8214 11994 8220 11996
rect 8276 11994 8300 11996
rect 8356 11994 8380 11996
rect 8436 11994 8460 11996
rect 8516 11994 8522 11996
rect 8276 11942 8278 11994
rect 8458 11942 8460 11994
rect 8214 11940 8220 11942
rect 8276 11940 8300 11942
rect 8356 11940 8380 11942
rect 8436 11940 8460 11942
rect 8516 11940 8522 11942
rect 8214 11931 8522 11940
rect 8588 11898 8616 12582
rect 9600 12458 9628 12974
rect 9876 12850 9904 13262
rect 10060 12918 10088 14962
rect 10336 14414 10364 15370
rect 10888 15162 10916 16526
rect 10980 16153 11008 17002
rect 10966 16144 11022 16153
rect 10966 16079 11022 16088
rect 11072 15706 11100 19314
rect 11440 19310 11468 19722
rect 11624 19446 11652 19790
rect 12256 19712 12308 19718
rect 12256 19654 12308 19660
rect 12268 19514 12296 19654
rect 12256 19508 12308 19514
rect 12256 19450 12308 19456
rect 11612 19440 11664 19446
rect 11612 19382 11664 19388
rect 11520 19372 11572 19378
rect 11520 19314 11572 19320
rect 11244 19304 11296 19310
rect 11244 19246 11296 19252
rect 11428 19304 11480 19310
rect 11428 19246 11480 19252
rect 11152 18964 11204 18970
rect 11152 18906 11204 18912
rect 11164 18698 11192 18906
rect 11256 18766 11284 19246
rect 11532 18766 11560 19314
rect 11624 19145 11652 19382
rect 12728 19378 12756 20198
rect 12992 19848 13044 19854
rect 12992 19790 13044 19796
rect 12072 19372 12124 19378
rect 11992 19332 12072 19360
rect 11610 19136 11666 19145
rect 11610 19071 11666 19080
rect 11888 18964 11940 18970
rect 11888 18906 11940 18912
rect 11702 18864 11758 18873
rect 11612 18828 11664 18834
rect 11702 18799 11758 18808
rect 11612 18770 11664 18776
rect 11244 18760 11296 18766
rect 11520 18760 11572 18766
rect 11244 18702 11296 18708
rect 11334 18728 11390 18737
rect 11152 18692 11204 18698
rect 11520 18702 11572 18708
rect 11334 18663 11390 18672
rect 11428 18692 11480 18698
rect 11152 18634 11204 18640
rect 11348 18272 11376 18663
rect 11428 18634 11480 18640
rect 11440 18601 11468 18634
rect 11426 18592 11482 18601
rect 11426 18527 11482 18536
rect 11426 18456 11482 18465
rect 11426 18391 11482 18400
rect 11440 18358 11468 18391
rect 11428 18352 11480 18358
rect 11428 18294 11480 18300
rect 11532 18290 11560 18702
rect 11624 18290 11652 18770
rect 11716 18766 11744 18799
rect 11704 18760 11756 18766
rect 11704 18702 11756 18708
rect 11256 18244 11376 18272
rect 11520 18284 11572 18290
rect 11152 18148 11204 18154
rect 11152 18090 11204 18096
rect 11164 17610 11192 18090
rect 11152 17604 11204 17610
rect 11152 17546 11204 17552
rect 11256 17202 11284 18244
rect 11520 18226 11572 18232
rect 11612 18284 11664 18290
rect 11612 18226 11664 18232
rect 11336 18148 11388 18154
rect 11336 18090 11388 18096
rect 11244 17196 11296 17202
rect 11244 17138 11296 17144
rect 11256 16561 11284 17138
rect 11348 17066 11376 18090
rect 11532 17882 11560 18226
rect 11610 17912 11666 17921
rect 11428 17876 11480 17882
rect 11428 17818 11480 17824
rect 11520 17876 11572 17882
rect 11900 17882 11928 18906
rect 11610 17847 11666 17856
rect 11888 17876 11940 17882
rect 11520 17818 11572 17824
rect 11440 17202 11468 17818
rect 11428 17196 11480 17202
rect 11428 17138 11480 17144
rect 11336 17060 11388 17066
rect 11336 17002 11388 17008
rect 11336 16584 11388 16590
rect 11242 16552 11298 16561
rect 11336 16526 11388 16532
rect 11242 16487 11298 16496
rect 11256 16454 11284 16487
rect 11244 16448 11296 16454
rect 11244 16390 11296 16396
rect 11348 16114 11376 16526
rect 11440 16114 11468 17138
rect 11532 16794 11560 17818
rect 11624 17066 11652 17847
rect 11888 17818 11940 17824
rect 11796 17536 11848 17542
rect 11794 17504 11796 17513
rect 11848 17504 11850 17513
rect 11794 17439 11850 17448
rect 11992 17252 12020 19332
rect 12072 19314 12124 19320
rect 12716 19372 12768 19378
rect 12716 19314 12768 19320
rect 12532 19168 12584 19174
rect 12584 19128 12664 19156
rect 12532 19110 12584 19116
rect 12214 19068 12522 19077
rect 12214 19066 12220 19068
rect 12276 19066 12300 19068
rect 12356 19066 12380 19068
rect 12436 19066 12460 19068
rect 12516 19066 12522 19068
rect 12276 19014 12278 19066
rect 12458 19014 12460 19066
rect 12214 19012 12220 19014
rect 12276 19012 12300 19014
rect 12356 19012 12380 19014
rect 12436 19012 12460 19014
rect 12516 19012 12522 19014
rect 12214 19003 12522 19012
rect 12636 18970 12664 19128
rect 12348 18964 12400 18970
rect 12348 18906 12400 18912
rect 12624 18964 12676 18970
rect 12624 18906 12676 18912
rect 12072 18896 12124 18902
rect 12070 18864 12072 18873
rect 12124 18864 12126 18873
rect 12070 18799 12126 18808
rect 12360 18766 12388 18906
rect 12438 18864 12494 18873
rect 12438 18799 12494 18808
rect 12452 18766 12480 18799
rect 12256 18760 12308 18766
rect 12256 18702 12308 18708
rect 12348 18760 12400 18766
rect 12348 18702 12400 18708
rect 12440 18760 12492 18766
rect 12624 18760 12676 18766
rect 12440 18702 12492 18708
rect 12622 18728 12624 18737
rect 12676 18728 12678 18737
rect 12268 18426 12296 18702
rect 12622 18663 12678 18672
rect 12346 18456 12402 18465
rect 12256 18420 12308 18426
rect 13004 18426 13032 19790
rect 13084 18896 13136 18902
rect 13084 18838 13136 18844
rect 12346 18391 12348 18400
rect 12256 18362 12308 18368
rect 12400 18391 12402 18400
rect 12992 18420 13044 18426
rect 12348 18362 12400 18368
rect 12992 18362 13044 18368
rect 12714 18320 12770 18329
rect 12072 18284 12124 18290
rect 12714 18255 12716 18264
rect 12072 18226 12124 18232
rect 12768 18255 12770 18264
rect 12808 18284 12860 18290
rect 12716 18226 12768 18232
rect 12860 18244 13032 18272
rect 12808 18226 12860 18232
rect 12084 18193 12112 18226
rect 12070 18184 12126 18193
rect 12070 18119 12126 18128
rect 12624 18148 12676 18154
rect 12624 18090 12676 18096
rect 12072 18080 12124 18086
rect 12072 18022 12124 18028
rect 12084 17864 12112 18022
rect 12214 17980 12522 17989
rect 12214 17978 12220 17980
rect 12276 17978 12300 17980
rect 12356 17978 12380 17980
rect 12436 17978 12460 17980
rect 12516 17978 12522 17980
rect 12276 17926 12278 17978
rect 12458 17926 12460 17978
rect 12214 17924 12220 17926
rect 12276 17924 12300 17926
rect 12356 17924 12380 17926
rect 12436 17924 12460 17926
rect 12516 17924 12522 17926
rect 12214 17915 12522 17924
rect 12084 17836 12296 17864
rect 12268 17542 12296 17836
rect 12164 17536 12216 17542
rect 12164 17478 12216 17484
rect 12256 17536 12308 17542
rect 12256 17478 12308 17484
rect 12176 17338 12204 17478
rect 12164 17332 12216 17338
rect 12164 17274 12216 17280
rect 11992 17224 12112 17252
rect 12084 17218 12112 17224
rect 12084 17190 12204 17218
rect 12636 17202 12664 18090
rect 13004 18086 13032 18244
rect 12716 18080 12768 18086
rect 12716 18022 12768 18028
rect 12992 18080 13044 18086
rect 12992 18022 13044 18028
rect 12728 17814 12756 18022
rect 13096 17882 13124 18838
rect 13188 18290 13216 21286
rect 13450 21200 13506 22000
rect 14556 21276 14608 21282
rect 14556 21218 14608 21224
rect 14280 21208 14332 21214
rect 13464 20058 13492 21200
rect 14280 21150 14332 21156
rect 14096 20800 14148 20806
rect 14096 20742 14148 20748
rect 13728 20460 13780 20466
rect 13728 20402 13780 20408
rect 13636 20392 13688 20398
rect 13636 20334 13688 20340
rect 13452 20052 13504 20058
rect 13452 19994 13504 20000
rect 13360 18760 13412 18766
rect 13360 18702 13412 18708
rect 13268 18692 13320 18698
rect 13268 18634 13320 18640
rect 13176 18284 13228 18290
rect 13176 18226 13228 18232
rect 12992 17876 13044 17882
rect 12992 17818 13044 17824
rect 13084 17876 13136 17882
rect 13084 17818 13136 17824
rect 12716 17808 12768 17814
rect 12716 17750 12768 17756
rect 12808 17808 12860 17814
rect 12808 17750 12860 17756
rect 12898 17776 12954 17785
rect 12716 17672 12768 17678
rect 12716 17614 12768 17620
rect 12728 17377 12756 17614
rect 12820 17542 12848 17750
rect 12898 17711 12954 17720
rect 12912 17542 12940 17711
rect 13004 17678 13032 17818
rect 13280 17814 13308 18634
rect 13372 18086 13400 18702
rect 13648 18630 13676 20334
rect 13740 19990 13768 20402
rect 13728 19984 13780 19990
rect 13728 19926 13780 19932
rect 13820 19780 13872 19786
rect 13820 19722 13872 19728
rect 13832 19514 13860 19722
rect 13820 19508 13872 19514
rect 13820 19450 13872 19456
rect 13818 18864 13874 18873
rect 13818 18799 13874 18808
rect 13832 18630 13860 18799
rect 14004 18760 14056 18766
rect 14004 18702 14056 18708
rect 13636 18624 13688 18630
rect 13636 18566 13688 18572
rect 13820 18624 13872 18630
rect 13872 18584 13952 18612
rect 13820 18566 13872 18572
rect 13556 18380 13768 18408
rect 13450 18320 13506 18329
rect 13450 18255 13506 18264
rect 13360 18080 13412 18086
rect 13360 18022 13412 18028
rect 13268 17808 13320 17814
rect 13268 17750 13320 17756
rect 12992 17672 13044 17678
rect 12992 17614 13044 17620
rect 13004 17542 13032 17614
rect 12808 17536 12860 17542
rect 12808 17478 12860 17484
rect 12900 17536 12952 17542
rect 12900 17478 12952 17484
rect 12992 17536 13044 17542
rect 12992 17478 13044 17484
rect 12714 17368 12770 17377
rect 12912 17338 12940 17478
rect 12714 17303 12770 17312
rect 12900 17332 12952 17338
rect 12900 17274 12952 17280
rect 12072 17128 12124 17134
rect 12072 17070 12124 17076
rect 11612 17060 11664 17066
rect 11612 17002 11664 17008
rect 11980 17060 12032 17066
rect 11980 17002 12032 17008
rect 11610 16824 11666 16833
rect 11520 16788 11572 16794
rect 11610 16759 11612 16768
rect 11520 16730 11572 16736
rect 11664 16759 11666 16768
rect 11888 16788 11940 16794
rect 11612 16730 11664 16736
rect 11888 16730 11940 16736
rect 11624 16658 11652 16730
rect 11612 16652 11664 16658
rect 11612 16594 11664 16600
rect 11520 16584 11572 16590
rect 11520 16526 11572 16532
rect 11336 16108 11388 16114
rect 11336 16050 11388 16056
rect 11428 16108 11480 16114
rect 11428 16050 11480 16056
rect 11152 16040 11204 16046
rect 11152 15982 11204 15988
rect 11060 15700 11112 15706
rect 11060 15642 11112 15648
rect 10968 15632 11020 15638
rect 11020 15580 11100 15586
rect 10968 15574 11100 15580
rect 10980 15558 11100 15574
rect 10876 15156 10928 15162
rect 10876 15098 10928 15104
rect 11072 14550 11100 15558
rect 11164 15484 11192 15982
rect 11348 15570 11376 16050
rect 11336 15564 11388 15570
rect 11336 15506 11388 15512
rect 11244 15496 11296 15502
rect 11164 15456 11244 15484
rect 11244 15438 11296 15444
rect 11152 15360 11204 15366
rect 11152 15302 11204 15308
rect 11164 15026 11192 15302
rect 11256 15026 11284 15438
rect 11348 15026 11376 15506
rect 11440 15162 11468 16050
rect 11532 15978 11560 16526
rect 11796 16448 11848 16454
rect 11900 16425 11928 16730
rect 11992 16726 12020 17002
rect 12084 16969 12112 17070
rect 12176 17066 12204 17190
rect 12624 17196 12676 17202
rect 12624 17138 12676 17144
rect 12808 17196 12860 17202
rect 12808 17138 12860 17144
rect 12900 17196 12952 17202
rect 12900 17138 12952 17144
rect 12164 17060 12216 17066
rect 12164 17002 12216 17008
rect 12070 16960 12126 16969
rect 12070 16895 12126 16904
rect 12214 16892 12522 16901
rect 12214 16890 12220 16892
rect 12276 16890 12300 16892
rect 12356 16890 12380 16892
rect 12436 16890 12460 16892
rect 12516 16890 12522 16892
rect 12276 16838 12278 16890
rect 12458 16838 12460 16890
rect 12214 16836 12220 16838
rect 12276 16836 12300 16838
rect 12356 16836 12380 16838
rect 12436 16836 12460 16838
rect 12516 16836 12522 16838
rect 12214 16827 12522 16836
rect 12820 16726 12848 17138
rect 11980 16720 12032 16726
rect 12256 16720 12308 16726
rect 11980 16662 12032 16668
rect 12070 16688 12126 16697
rect 12256 16662 12308 16668
rect 12624 16720 12676 16726
rect 12624 16662 12676 16668
rect 12808 16720 12860 16726
rect 12808 16662 12860 16668
rect 12070 16623 12126 16632
rect 12084 16522 12112 16623
rect 12164 16584 12216 16590
rect 12162 16552 12164 16561
rect 12216 16552 12218 16561
rect 12072 16516 12124 16522
rect 12268 16522 12296 16662
rect 12532 16584 12584 16590
rect 12532 16526 12584 16532
rect 12162 16487 12218 16496
rect 12256 16516 12308 16522
rect 12072 16458 12124 16464
rect 12256 16458 12308 16464
rect 11796 16390 11848 16396
rect 11886 16416 11942 16425
rect 11610 16280 11666 16289
rect 11808 16250 11836 16390
rect 11886 16351 11942 16360
rect 11610 16215 11612 16224
rect 11664 16215 11666 16224
rect 11796 16244 11848 16250
rect 11612 16186 11664 16192
rect 11796 16186 11848 16192
rect 11980 16176 12032 16182
rect 11980 16118 12032 16124
rect 11520 15972 11572 15978
rect 11520 15914 11572 15920
rect 11704 15904 11756 15910
rect 11704 15846 11756 15852
rect 11716 15502 11744 15846
rect 11704 15496 11756 15502
rect 11704 15438 11756 15444
rect 11888 15496 11940 15502
rect 11888 15438 11940 15444
rect 11428 15156 11480 15162
rect 11428 15098 11480 15104
rect 11152 15020 11204 15026
rect 11152 14962 11204 14968
rect 11244 15020 11296 15026
rect 11244 14962 11296 14968
rect 11336 15020 11388 15026
rect 11336 14962 11388 14968
rect 11900 14550 11928 15438
rect 11992 15162 12020 16118
rect 12084 16046 12112 16458
rect 12440 16448 12492 16454
rect 12440 16390 12492 16396
rect 12452 16114 12480 16390
rect 12544 16182 12572 16526
rect 12532 16176 12584 16182
rect 12532 16118 12584 16124
rect 12440 16108 12492 16114
rect 12440 16050 12492 16056
rect 12072 16040 12124 16046
rect 12072 15982 12124 15988
rect 12214 15804 12522 15813
rect 12214 15802 12220 15804
rect 12276 15802 12300 15804
rect 12356 15802 12380 15804
rect 12436 15802 12460 15804
rect 12516 15802 12522 15804
rect 12276 15750 12278 15802
rect 12458 15750 12460 15802
rect 12214 15748 12220 15750
rect 12276 15748 12300 15750
rect 12356 15748 12380 15750
rect 12436 15748 12460 15750
rect 12516 15748 12522 15750
rect 12214 15739 12522 15748
rect 12440 15632 12492 15638
rect 12636 15586 12664 16662
rect 12808 16584 12860 16590
rect 12728 16544 12808 16572
rect 12728 16114 12756 16544
rect 12912 16572 12940 17138
rect 13004 16726 13032 17478
rect 13268 17128 13320 17134
rect 13268 17070 13320 17076
rect 12992 16720 13044 16726
rect 12992 16662 13044 16668
rect 13176 16584 13228 16590
rect 12860 16544 13176 16572
rect 12808 16526 12860 16532
rect 13176 16526 13228 16532
rect 13280 16250 13308 17070
rect 13372 16250 13400 18022
rect 13464 17678 13492 18255
rect 13452 17672 13504 17678
rect 13452 17614 13504 17620
rect 13464 17202 13492 17614
rect 13452 17196 13504 17202
rect 13452 17138 13504 17144
rect 13556 17105 13584 18380
rect 13740 18290 13768 18380
rect 13636 18284 13688 18290
rect 13636 18226 13688 18232
rect 13728 18284 13780 18290
rect 13728 18226 13780 18232
rect 13820 18284 13872 18290
rect 13820 18226 13872 18232
rect 13648 17678 13676 18226
rect 13832 17746 13860 18226
rect 13820 17740 13872 17746
rect 13820 17682 13872 17688
rect 13636 17672 13688 17678
rect 13636 17614 13688 17620
rect 13818 17640 13874 17649
rect 13648 17513 13676 17614
rect 13818 17575 13820 17584
rect 13872 17575 13874 17584
rect 13820 17546 13872 17552
rect 13924 17542 13952 18584
rect 13912 17536 13964 17542
rect 13634 17504 13690 17513
rect 13912 17478 13964 17484
rect 13634 17439 13690 17448
rect 14016 17338 14044 18702
rect 14108 17338 14136 20742
rect 14188 20324 14240 20330
rect 14188 20266 14240 20272
rect 14200 20058 14228 20266
rect 14188 20052 14240 20058
rect 14188 19994 14240 20000
rect 14188 19780 14240 19786
rect 14188 19722 14240 19728
rect 14200 19378 14228 19722
rect 14188 19372 14240 19378
rect 14188 19314 14240 19320
rect 14200 18970 14228 19314
rect 14188 18964 14240 18970
rect 14188 18906 14240 18912
rect 14292 18358 14320 21150
rect 14568 18766 14596 21218
rect 15474 21200 15530 22000
rect 17498 21298 17554 22000
rect 17328 21270 17554 21298
rect 15292 20936 15344 20942
rect 15292 20878 15344 20884
rect 14648 20868 14700 20874
rect 14648 20810 14700 20816
rect 14556 18760 14608 18766
rect 14556 18702 14608 18708
rect 14280 18352 14332 18358
rect 14280 18294 14332 18300
rect 14556 18284 14608 18290
rect 14556 18226 14608 18232
rect 14372 18216 14424 18222
rect 14372 18158 14424 18164
rect 14384 17678 14412 18158
rect 14568 18154 14596 18226
rect 14556 18148 14608 18154
rect 14556 18090 14608 18096
rect 14660 17678 14688 20810
rect 15016 20256 15068 20262
rect 15016 20198 15068 20204
rect 15200 20256 15252 20262
rect 15200 20198 15252 20204
rect 15028 19990 15056 20198
rect 15016 19984 15068 19990
rect 15016 19926 15068 19932
rect 15028 19378 15056 19926
rect 15212 19922 15240 20198
rect 15200 19916 15252 19922
rect 15200 19858 15252 19864
rect 15016 19372 15068 19378
rect 15016 19314 15068 19320
rect 15200 18692 15252 18698
rect 15200 18634 15252 18640
rect 15212 18426 15240 18634
rect 15200 18420 15252 18426
rect 15200 18362 15252 18368
rect 15200 18284 15252 18290
rect 15304 18272 15332 20878
rect 15488 20618 15516 21200
rect 15568 21004 15620 21010
rect 15568 20946 15620 20952
rect 15396 20590 15516 20618
rect 15396 20058 15424 20590
rect 15476 20460 15528 20466
rect 15476 20402 15528 20408
rect 15488 20058 15516 20402
rect 15384 20052 15436 20058
rect 15384 19994 15436 20000
rect 15476 20052 15528 20058
rect 15476 19994 15528 20000
rect 15476 19780 15528 19786
rect 15476 19722 15528 19728
rect 15488 19446 15516 19722
rect 15476 19440 15528 19446
rect 15476 19382 15528 19388
rect 15384 19304 15436 19310
rect 15384 19246 15436 19252
rect 15252 18244 15332 18272
rect 15200 18226 15252 18232
rect 15396 18222 15424 19246
rect 15474 18592 15530 18601
rect 15474 18527 15530 18536
rect 15488 18426 15516 18527
rect 15476 18420 15528 18426
rect 15476 18362 15528 18368
rect 15476 18284 15528 18290
rect 15476 18226 15528 18232
rect 15384 18216 15436 18222
rect 15384 18158 15436 18164
rect 15488 17814 15516 18226
rect 15580 17882 15608 20946
rect 16214 20700 16522 20709
rect 16214 20698 16220 20700
rect 16276 20698 16300 20700
rect 16356 20698 16380 20700
rect 16436 20698 16460 20700
rect 16516 20698 16522 20700
rect 16276 20646 16278 20698
rect 16458 20646 16460 20698
rect 16214 20644 16220 20646
rect 16276 20644 16300 20646
rect 16356 20644 16380 20646
rect 16436 20644 16460 20646
rect 16516 20644 16522 20646
rect 16214 20635 16522 20644
rect 16304 20596 16356 20602
rect 16304 20538 16356 20544
rect 15660 20392 15712 20398
rect 15660 20334 15712 20340
rect 15752 20392 15804 20398
rect 15752 20334 15804 20340
rect 15672 19922 15700 20334
rect 15660 19916 15712 19922
rect 15660 19858 15712 19864
rect 15764 19718 15792 20334
rect 16316 20058 16344 20538
rect 17224 20324 17276 20330
rect 17224 20266 17276 20272
rect 17236 20058 17264 20266
rect 16304 20052 16356 20058
rect 16304 19994 16356 20000
rect 17224 20052 17276 20058
rect 17224 19994 17276 20000
rect 16672 19984 16724 19990
rect 16672 19926 16724 19932
rect 16684 19825 16712 19926
rect 16670 19816 16726 19825
rect 16580 19780 16632 19786
rect 16670 19751 16726 19760
rect 16580 19722 16632 19728
rect 15752 19712 15804 19718
rect 15752 19654 15804 19660
rect 16214 19612 16522 19621
rect 16214 19610 16220 19612
rect 16276 19610 16300 19612
rect 16356 19610 16380 19612
rect 16436 19610 16460 19612
rect 16516 19610 16522 19612
rect 16276 19558 16278 19610
rect 16458 19558 16460 19610
rect 16214 19556 16220 19558
rect 16276 19556 16300 19558
rect 16356 19556 16380 19558
rect 16436 19556 16460 19558
rect 16516 19556 16522 19558
rect 16214 19547 16522 19556
rect 16592 19514 16620 19722
rect 16764 19712 16816 19718
rect 16764 19654 16816 19660
rect 16580 19508 16632 19514
rect 16580 19450 16632 19456
rect 16776 19446 16804 19654
rect 16764 19440 16816 19446
rect 16764 19382 16816 19388
rect 16028 19304 16080 19310
rect 16396 19304 16448 19310
rect 16080 19252 16396 19258
rect 16028 19246 16448 19252
rect 16040 19230 16436 19246
rect 16764 19236 16816 19242
rect 16764 19178 16816 19184
rect 16776 18766 16804 19178
rect 16764 18760 16816 18766
rect 16764 18702 16816 18708
rect 16948 18624 17000 18630
rect 16948 18566 17000 18572
rect 17224 18624 17276 18630
rect 17224 18566 17276 18572
rect 16214 18524 16522 18533
rect 16214 18522 16220 18524
rect 16276 18522 16300 18524
rect 16356 18522 16380 18524
rect 16436 18522 16460 18524
rect 16516 18522 16522 18524
rect 16276 18470 16278 18522
rect 16458 18470 16460 18522
rect 16214 18468 16220 18470
rect 16276 18468 16300 18470
rect 16356 18468 16380 18470
rect 16436 18468 16460 18470
rect 16516 18468 16522 18470
rect 16214 18459 16522 18468
rect 16960 18358 16988 18566
rect 16948 18352 17000 18358
rect 16948 18294 17000 18300
rect 16028 18216 16080 18222
rect 16028 18158 16080 18164
rect 16040 17882 16068 18158
rect 15568 17876 15620 17882
rect 15568 17818 15620 17824
rect 16028 17876 16080 17882
rect 16028 17818 16080 17824
rect 17236 17814 17264 18566
rect 15476 17808 15528 17814
rect 15476 17750 15528 17756
rect 17224 17808 17276 17814
rect 17224 17750 17276 17756
rect 14372 17672 14424 17678
rect 14372 17614 14424 17620
rect 14648 17672 14700 17678
rect 14648 17614 14700 17620
rect 15568 17672 15620 17678
rect 15568 17614 15620 17620
rect 16028 17672 16080 17678
rect 16028 17614 16080 17620
rect 14464 17604 14516 17610
rect 14464 17546 14516 17552
rect 14280 17536 14332 17542
rect 14280 17478 14332 17484
rect 14004 17332 14056 17338
rect 14004 17274 14056 17280
rect 14096 17332 14148 17338
rect 14096 17274 14148 17280
rect 14292 17270 14320 17478
rect 14280 17264 14332 17270
rect 14280 17206 14332 17212
rect 13728 17196 13780 17202
rect 13728 17138 13780 17144
rect 14188 17196 14240 17202
rect 14188 17138 14240 17144
rect 13542 17096 13598 17105
rect 13542 17031 13598 17040
rect 13556 16658 13584 17031
rect 13544 16652 13596 16658
rect 13544 16594 13596 16600
rect 13740 16590 13768 17138
rect 13728 16584 13780 16590
rect 13728 16526 13780 16532
rect 12992 16244 13044 16250
rect 12992 16186 13044 16192
rect 13268 16244 13320 16250
rect 13268 16186 13320 16192
rect 13360 16244 13412 16250
rect 13360 16186 13412 16192
rect 12716 16108 12768 16114
rect 12716 16050 12768 16056
rect 12808 16108 12860 16114
rect 12808 16050 12860 16056
rect 12492 15580 12664 15586
rect 12440 15574 12664 15580
rect 12452 15558 12664 15574
rect 12728 15502 12756 16050
rect 12716 15496 12768 15502
rect 12716 15438 12768 15444
rect 12820 15366 12848 16050
rect 12900 16040 12952 16046
rect 12900 15982 12952 15988
rect 12912 15706 12940 15982
rect 13004 15910 13032 16186
rect 13740 16046 13768 16526
rect 14200 16250 14228 17138
rect 14476 16697 14504 17546
rect 14832 17536 14884 17542
rect 14832 17478 14884 17484
rect 14844 17270 14872 17478
rect 14832 17264 14884 17270
rect 14832 17206 14884 17212
rect 15382 17232 15438 17241
rect 15382 17167 15438 17176
rect 14556 16992 14608 16998
rect 14556 16934 14608 16940
rect 14462 16688 14518 16697
rect 14462 16623 14518 16632
rect 14188 16244 14240 16250
rect 14188 16186 14240 16192
rect 14568 16182 14596 16934
rect 14924 16720 14976 16726
rect 14976 16680 15148 16708
rect 14924 16662 14976 16668
rect 15120 16590 15148 16680
rect 15108 16584 15160 16590
rect 15108 16526 15160 16532
rect 15120 16250 15148 16526
rect 15396 16522 15424 17167
rect 15384 16516 15436 16522
rect 15384 16458 15436 16464
rect 15108 16244 15160 16250
rect 15108 16186 15160 16192
rect 14556 16176 14608 16182
rect 14556 16118 14608 16124
rect 13728 16040 13780 16046
rect 13728 15982 13780 15988
rect 12992 15904 13044 15910
rect 12992 15846 13044 15852
rect 12900 15700 12952 15706
rect 12900 15642 12952 15648
rect 13084 15632 13136 15638
rect 13084 15574 13136 15580
rect 13096 15434 13124 15574
rect 13740 15570 13768 15982
rect 14568 15570 14596 16118
rect 15108 16108 15160 16114
rect 15108 16050 15160 16056
rect 13728 15564 13780 15570
rect 13728 15506 13780 15512
rect 14556 15564 14608 15570
rect 14556 15506 14608 15512
rect 13636 15496 13688 15502
rect 13636 15438 13688 15444
rect 13084 15428 13136 15434
rect 13084 15370 13136 15376
rect 13176 15428 13228 15434
rect 13176 15370 13228 15376
rect 12808 15360 12860 15366
rect 12808 15302 12860 15308
rect 12820 15162 12848 15302
rect 11980 15156 12032 15162
rect 11980 15098 12032 15104
rect 12808 15156 12860 15162
rect 12808 15098 12860 15104
rect 12072 15020 12124 15026
rect 12072 14962 12124 14968
rect 11060 14544 11112 14550
rect 11060 14486 11112 14492
rect 11888 14544 11940 14550
rect 11888 14486 11940 14492
rect 10784 14476 10836 14482
rect 10784 14418 10836 14424
rect 10324 14408 10376 14414
rect 10324 14350 10376 14356
rect 10796 14346 10824 14418
rect 10784 14340 10836 14346
rect 10784 14282 10836 14288
rect 10508 13728 10560 13734
rect 10508 13670 10560 13676
rect 10416 13388 10468 13394
rect 10416 13330 10468 13336
rect 10048 12912 10100 12918
rect 10048 12854 10100 12860
rect 9680 12844 9732 12850
rect 9680 12786 9732 12792
rect 9864 12844 9916 12850
rect 9864 12786 9916 12792
rect 9692 12594 9720 12786
rect 9692 12566 9812 12594
rect 9600 12430 9720 12458
rect 9692 12238 9720 12430
rect 9784 12374 9812 12566
rect 9772 12368 9824 12374
rect 9772 12310 9824 12316
rect 9680 12232 9732 12238
rect 9680 12174 9732 12180
rect 9772 12096 9824 12102
rect 9772 12038 9824 12044
rect 8576 11892 8628 11898
rect 8576 11834 8628 11840
rect 9784 11830 9812 12038
rect 10060 11898 10088 12854
rect 10140 12368 10192 12374
rect 10140 12310 10192 12316
rect 10048 11892 10100 11898
rect 10048 11834 10100 11840
rect 9772 11824 9824 11830
rect 9772 11766 9824 11772
rect 7840 11756 7892 11762
rect 7840 11698 7892 11704
rect 7852 11286 7880 11698
rect 9956 11552 10008 11558
rect 9956 11494 10008 11500
rect 9968 11354 9996 11494
rect 9956 11348 10008 11354
rect 9956 11290 10008 11296
rect 7748 11280 7800 11286
rect 7748 11222 7800 11228
rect 7840 11280 7892 11286
rect 7840 11222 7892 11228
rect 7380 11212 7432 11218
rect 7380 11154 7432 11160
rect 6828 11144 6880 11150
rect 6828 11086 6880 11092
rect 7012 11144 7064 11150
rect 7012 11086 7064 11092
rect 7392 10810 7420 11154
rect 6920 10804 6972 10810
rect 6920 10746 6972 10752
rect 7380 10804 7432 10810
rect 7380 10746 7432 10752
rect 6932 10266 6960 10746
rect 6920 10260 6972 10266
rect 6920 10202 6972 10208
rect 6920 10056 6972 10062
rect 6656 9710 6776 9738
rect 6840 10016 6920 10044
rect 6552 9648 6604 9654
rect 6552 9590 6604 9596
rect 6564 9178 6592 9590
rect 6552 9172 6604 9178
rect 6552 9114 6604 9120
rect 6368 8084 6420 8090
rect 6368 8026 6420 8032
rect 6368 7880 6420 7886
rect 6368 7822 6420 7828
rect 6000 7812 6052 7818
rect 6000 7754 6052 7760
rect 6012 7002 6040 7754
rect 6092 7540 6144 7546
rect 6092 7482 6144 7488
rect 6000 6996 6052 7002
rect 6000 6938 6052 6944
rect 6104 6798 6132 7482
rect 6276 7472 6328 7478
rect 6380 7460 6408 7822
rect 6656 7562 6684 9710
rect 6736 9580 6788 9586
rect 6736 9522 6788 9528
rect 6748 9178 6776 9522
rect 6840 9518 6868 10016
rect 6920 9998 6972 10004
rect 7564 10056 7616 10062
rect 7564 9998 7616 10004
rect 7196 9580 7248 9586
rect 7196 9522 7248 9528
rect 6828 9512 6880 9518
rect 6828 9454 6880 9460
rect 6736 9172 6788 9178
rect 6736 9114 6788 9120
rect 7104 8968 7156 8974
rect 7104 8910 7156 8916
rect 7116 8634 7144 8910
rect 7104 8628 7156 8634
rect 7104 8570 7156 8576
rect 7116 8498 7144 8570
rect 7208 8498 7236 9522
rect 7576 9382 7604 9998
rect 7760 9518 7788 11222
rect 7852 10674 7880 11222
rect 7932 11144 7984 11150
rect 7932 11086 7984 11092
rect 9036 11144 9088 11150
rect 9036 11086 9088 11092
rect 7840 10668 7892 10674
rect 7840 10610 7892 10616
rect 7852 9654 7880 10610
rect 7944 10266 7972 11086
rect 8116 11008 8168 11014
rect 8116 10950 8168 10956
rect 8024 10804 8076 10810
rect 8024 10746 8076 10752
rect 7932 10260 7984 10266
rect 7932 10202 7984 10208
rect 7932 10056 7984 10062
rect 7932 9998 7984 10004
rect 7840 9648 7892 9654
rect 7840 9590 7892 9596
rect 7748 9512 7800 9518
rect 7748 9454 7800 9460
rect 7564 9376 7616 9382
rect 7564 9318 7616 9324
rect 7852 9042 7880 9590
rect 7840 9036 7892 9042
rect 7840 8978 7892 8984
rect 7288 8832 7340 8838
rect 7288 8774 7340 8780
rect 7104 8492 7156 8498
rect 7104 8434 7156 8440
rect 7196 8492 7248 8498
rect 7196 8434 7248 8440
rect 6328 7432 6408 7460
rect 6276 7414 6328 7420
rect 6092 6792 6144 6798
rect 6092 6734 6144 6740
rect 6092 6656 6144 6662
rect 6092 6598 6144 6604
rect 6104 5710 6132 6598
rect 6380 6458 6408 7432
rect 6564 7534 6684 7562
rect 7104 7540 7156 7546
rect 6368 6452 6420 6458
rect 6368 6394 6420 6400
rect 6092 5704 6144 5710
rect 6092 5646 6144 5652
rect 6000 5636 6052 5642
rect 6000 5578 6052 5584
rect 5908 5568 5960 5574
rect 5908 5510 5960 5516
rect 6012 5234 6040 5578
rect 6000 5228 6052 5234
rect 6000 5170 6052 5176
rect 5264 4752 5316 4758
rect 5264 4694 5316 4700
rect 5540 4752 5592 4758
rect 5540 4694 5592 4700
rect 6276 4004 6328 4010
rect 6276 3946 6328 3952
rect 6184 3664 6236 3670
rect 6184 3606 6236 3612
rect 6196 3534 6224 3606
rect 6288 3534 6316 3946
rect 6184 3528 6236 3534
rect 6184 3470 6236 3476
rect 6276 3528 6328 3534
rect 6276 3470 6328 3476
rect 5906 3360 5962 3369
rect 5906 3295 5962 3304
rect 5172 3188 5224 3194
rect 5172 3130 5224 3136
rect 5920 3058 5948 3295
rect 5908 3052 5960 3058
rect 5908 2994 5960 3000
rect 5632 2984 5684 2990
rect 5632 2926 5684 2932
rect 5644 2106 5672 2926
rect 5632 2100 5684 2106
rect 5632 2042 5684 2048
rect 5920 1970 5948 2994
rect 6000 2984 6052 2990
rect 6000 2926 6052 2932
rect 6012 2446 6040 2926
rect 6564 2774 6592 7534
rect 7104 7482 7156 7488
rect 6644 7404 6696 7410
rect 6644 7346 6696 7352
rect 7012 7404 7064 7410
rect 7012 7346 7064 7352
rect 6656 6934 6684 7346
rect 6644 6928 6696 6934
rect 6644 6870 6696 6876
rect 7024 6458 7052 7346
rect 7116 7002 7144 7482
rect 7208 7342 7236 8434
rect 7196 7336 7248 7342
rect 7196 7278 7248 7284
rect 7104 6996 7156 7002
rect 7104 6938 7156 6944
rect 7116 6662 7144 6938
rect 7104 6656 7156 6662
rect 7104 6598 7156 6604
rect 7012 6452 7064 6458
rect 7012 6394 7064 6400
rect 7104 6316 7156 6322
rect 7104 6258 7156 6264
rect 7116 5914 7144 6258
rect 7104 5908 7156 5914
rect 7104 5850 7156 5856
rect 6920 5840 6972 5846
rect 7300 5794 7328 8774
rect 7380 8560 7432 8566
rect 7380 8502 7432 8508
rect 7392 6866 7420 8502
rect 7748 7744 7800 7750
rect 7748 7686 7800 7692
rect 7472 7200 7524 7206
rect 7472 7142 7524 7148
rect 7484 6866 7512 7142
rect 7380 6860 7432 6866
rect 7380 6802 7432 6808
rect 7472 6860 7524 6866
rect 7472 6802 7524 6808
rect 7760 6798 7788 7686
rect 7748 6792 7800 6798
rect 7748 6734 7800 6740
rect 7840 6384 7892 6390
rect 7944 6372 7972 9998
rect 8036 8974 8064 10746
rect 8128 10742 8156 10950
rect 8214 10908 8522 10917
rect 8214 10906 8220 10908
rect 8276 10906 8300 10908
rect 8356 10906 8380 10908
rect 8436 10906 8460 10908
rect 8516 10906 8522 10908
rect 8276 10854 8278 10906
rect 8458 10854 8460 10906
rect 8214 10852 8220 10854
rect 8276 10852 8300 10854
rect 8356 10852 8380 10854
rect 8436 10852 8460 10854
rect 8516 10852 8522 10854
rect 8214 10843 8522 10852
rect 8116 10736 8168 10742
rect 8116 10678 8168 10684
rect 9048 10266 9076 11086
rect 9312 11076 9364 11082
rect 9312 11018 9364 11024
rect 9036 10260 9088 10266
rect 9036 10202 9088 10208
rect 9220 10260 9272 10266
rect 9220 10202 9272 10208
rect 8760 9988 8812 9994
rect 8760 9930 8812 9936
rect 8214 9820 8522 9829
rect 8214 9818 8220 9820
rect 8276 9818 8300 9820
rect 8356 9818 8380 9820
rect 8436 9818 8460 9820
rect 8516 9818 8522 9820
rect 8276 9766 8278 9818
rect 8458 9766 8460 9818
rect 8214 9764 8220 9766
rect 8276 9764 8300 9766
rect 8356 9764 8380 9766
rect 8436 9764 8460 9766
rect 8516 9764 8522 9766
rect 8214 9755 8522 9764
rect 8024 8968 8076 8974
rect 8024 8910 8076 8916
rect 8214 8732 8522 8741
rect 8214 8730 8220 8732
rect 8276 8730 8300 8732
rect 8356 8730 8380 8732
rect 8436 8730 8460 8732
rect 8516 8730 8522 8732
rect 8276 8678 8278 8730
rect 8458 8678 8460 8730
rect 8214 8676 8220 8678
rect 8276 8676 8300 8678
rect 8356 8676 8380 8678
rect 8436 8676 8460 8678
rect 8516 8676 8522 8678
rect 8214 8667 8522 8676
rect 8300 8628 8352 8634
rect 8300 8570 8352 8576
rect 8312 7886 8340 8570
rect 8772 8362 8800 9930
rect 9232 9926 9260 10202
rect 9220 9920 9272 9926
rect 9220 9862 9272 9868
rect 9232 9722 9260 9862
rect 9220 9716 9272 9722
rect 9220 9658 9272 9664
rect 9324 9654 9352 11018
rect 9864 11008 9916 11014
rect 9864 10950 9916 10956
rect 10048 11008 10100 11014
rect 10048 10950 10100 10956
rect 9876 10674 9904 10950
rect 10060 10674 10088 10950
rect 9864 10668 9916 10674
rect 9864 10610 9916 10616
rect 10048 10668 10100 10674
rect 10048 10610 10100 10616
rect 9496 10532 9548 10538
rect 9496 10474 9548 10480
rect 9404 10464 9456 10470
rect 9404 10406 9456 10412
rect 9312 9648 9364 9654
rect 9312 9590 9364 9596
rect 9312 8424 9364 8430
rect 9312 8366 9364 8372
rect 8760 8356 8812 8362
rect 8760 8298 8812 8304
rect 8576 7948 8628 7954
rect 8576 7890 8628 7896
rect 8116 7880 8168 7886
rect 8116 7822 8168 7828
rect 8300 7880 8352 7886
rect 8300 7822 8352 7828
rect 8024 7744 8076 7750
rect 8024 7686 8076 7692
rect 8036 7478 8064 7686
rect 8024 7472 8076 7478
rect 8024 7414 8076 7420
rect 8128 7290 8156 7822
rect 8214 7644 8522 7653
rect 8214 7642 8220 7644
rect 8276 7642 8300 7644
rect 8356 7642 8380 7644
rect 8436 7642 8460 7644
rect 8516 7642 8522 7644
rect 8276 7590 8278 7642
rect 8458 7590 8460 7642
rect 8214 7588 8220 7590
rect 8276 7588 8300 7590
rect 8356 7588 8380 7590
rect 8436 7588 8460 7590
rect 8516 7588 8522 7590
rect 8214 7579 8522 7588
rect 8036 7262 8156 7290
rect 8036 6798 8064 7262
rect 8588 6798 8616 7890
rect 8668 7880 8720 7886
rect 8668 7822 8720 7828
rect 8680 6866 8708 7822
rect 8772 6934 8800 8298
rect 8944 7744 8996 7750
rect 8944 7686 8996 7692
rect 8760 6928 8812 6934
rect 8760 6870 8812 6876
rect 8668 6860 8720 6866
rect 8668 6802 8720 6808
rect 8024 6792 8076 6798
rect 8024 6734 8076 6740
rect 8576 6792 8628 6798
rect 8772 6746 8800 6870
rect 8576 6734 8628 6740
rect 7892 6344 7972 6372
rect 8036 6372 8064 6734
rect 8680 6730 8800 6746
rect 8668 6724 8800 6730
rect 8720 6718 8800 6724
rect 8668 6666 8720 6672
rect 8576 6656 8628 6662
rect 8576 6598 8628 6604
rect 8852 6656 8904 6662
rect 8852 6598 8904 6604
rect 8214 6556 8522 6565
rect 8214 6554 8220 6556
rect 8276 6554 8300 6556
rect 8356 6554 8380 6556
rect 8436 6554 8460 6556
rect 8516 6554 8522 6556
rect 8276 6502 8278 6554
rect 8458 6502 8460 6554
rect 8214 6500 8220 6502
rect 8276 6500 8300 6502
rect 8356 6500 8380 6502
rect 8436 6500 8460 6502
rect 8516 6500 8522 6502
rect 8214 6491 8522 6500
rect 8208 6384 8260 6390
rect 8036 6344 8208 6372
rect 7840 6326 7892 6332
rect 7656 6112 7708 6118
rect 7656 6054 7708 6060
rect 7748 6112 7800 6118
rect 7748 6054 7800 6060
rect 6920 5782 6972 5788
rect 6932 5302 6960 5782
rect 7208 5766 7328 5794
rect 7012 5636 7064 5642
rect 7012 5578 7064 5584
rect 7104 5636 7156 5642
rect 7104 5578 7156 5584
rect 7024 5370 7052 5578
rect 7012 5364 7064 5370
rect 7012 5306 7064 5312
rect 6920 5296 6972 5302
rect 6920 5238 6972 5244
rect 7116 5098 7144 5578
rect 7104 5092 7156 5098
rect 7104 5034 7156 5040
rect 7012 5024 7064 5030
rect 7208 4978 7236 5766
rect 7380 5704 7432 5710
rect 7380 5646 7432 5652
rect 7392 5166 7420 5646
rect 7564 5636 7616 5642
rect 7564 5578 7616 5584
rect 7576 5234 7604 5578
rect 7668 5574 7696 6054
rect 7760 5574 7788 6054
rect 7852 5710 7880 6326
rect 7840 5704 7892 5710
rect 7840 5646 7892 5652
rect 7656 5568 7708 5574
rect 7656 5510 7708 5516
rect 7748 5568 7800 5574
rect 7748 5510 7800 5516
rect 7852 5370 7880 5646
rect 8036 5642 8064 6344
rect 8208 6326 8260 6332
rect 8300 6316 8352 6322
rect 8300 6258 8352 6264
rect 8208 6112 8260 6118
rect 8208 6054 8260 6060
rect 8220 5710 8248 6054
rect 8312 5778 8340 6258
rect 8588 6254 8616 6598
rect 8864 6322 8892 6598
rect 8956 6390 8984 7686
rect 9036 7336 9088 7342
rect 9036 7278 9088 7284
rect 8944 6384 8996 6390
rect 8944 6326 8996 6332
rect 8760 6316 8812 6322
rect 8760 6258 8812 6264
rect 8852 6316 8904 6322
rect 8852 6258 8904 6264
rect 8576 6248 8628 6254
rect 8576 6190 8628 6196
rect 8772 6186 8800 6258
rect 8760 6180 8812 6186
rect 8760 6122 8812 6128
rect 8668 6112 8720 6118
rect 8668 6054 8720 6060
rect 8300 5772 8352 5778
rect 8300 5714 8352 5720
rect 8208 5704 8260 5710
rect 8208 5646 8260 5652
rect 8024 5636 8076 5642
rect 8024 5578 8076 5584
rect 8214 5468 8522 5477
rect 8214 5466 8220 5468
rect 8276 5466 8300 5468
rect 8356 5466 8380 5468
rect 8436 5466 8460 5468
rect 8516 5466 8522 5468
rect 8276 5414 8278 5466
rect 8458 5414 8460 5466
rect 8214 5412 8220 5414
rect 8276 5412 8300 5414
rect 8356 5412 8380 5414
rect 8436 5412 8460 5414
rect 8516 5412 8522 5414
rect 8214 5403 8522 5412
rect 7656 5364 7708 5370
rect 7656 5306 7708 5312
rect 7840 5364 7892 5370
rect 7840 5306 7892 5312
rect 7564 5228 7616 5234
rect 7564 5170 7616 5176
rect 7380 5160 7432 5166
rect 7380 5102 7432 5108
rect 7012 4966 7064 4972
rect 7024 4622 7052 4966
rect 7116 4950 7236 4978
rect 7012 4616 7064 4622
rect 7012 4558 7064 4564
rect 7116 4078 7144 4950
rect 7196 4616 7248 4622
rect 7196 4558 7248 4564
rect 7208 4486 7236 4558
rect 7196 4480 7248 4486
rect 7196 4422 7248 4428
rect 7208 4282 7236 4422
rect 7196 4276 7248 4282
rect 7196 4218 7248 4224
rect 6644 4072 6696 4078
rect 6644 4014 6696 4020
rect 7104 4072 7156 4078
rect 7104 4014 7156 4020
rect 6656 3738 6684 4014
rect 6644 3732 6696 3738
rect 6644 3674 6696 3680
rect 6736 3120 6788 3126
rect 6736 3062 6788 3068
rect 6564 2746 6684 2774
rect 6000 2440 6052 2446
rect 6000 2382 6052 2388
rect 6012 1970 6040 2382
rect 6460 2372 6512 2378
rect 6460 2314 6512 2320
rect 6276 2304 6328 2310
rect 6276 2246 6328 2252
rect 5908 1964 5960 1970
rect 5908 1906 5960 1912
rect 6000 1964 6052 1970
rect 6000 1906 6052 1912
rect 6288 1902 6316 2246
rect 6276 1896 6328 1902
rect 6276 1838 6328 1844
rect 6472 1834 6500 2314
rect 5080 1828 5132 1834
rect 5080 1770 5132 1776
rect 6460 1828 6512 1834
rect 6460 1770 6512 1776
rect 4988 1556 5040 1562
rect 4988 1498 5040 1504
rect 5092 1358 5120 1770
rect 2872 1352 2924 1358
rect 846 1320 902 1329
rect 2872 1294 2924 1300
rect 4896 1352 4948 1358
rect 4896 1294 4948 1300
rect 5080 1352 5132 1358
rect 5080 1294 5132 1300
rect 846 1255 902 1264
rect 6656 1170 6684 2746
rect 6748 2378 6776 3062
rect 7116 2774 7144 4014
rect 7392 3738 7420 5102
rect 7668 4826 7696 5306
rect 7932 5228 7984 5234
rect 7932 5170 7984 5176
rect 7944 4826 7972 5170
rect 8484 5024 8536 5030
rect 8484 4966 8536 4972
rect 7656 4820 7708 4826
rect 7656 4762 7708 4768
rect 7932 4820 7984 4826
rect 7932 4762 7984 4768
rect 8496 4622 8524 4966
rect 8484 4616 8536 4622
rect 8484 4558 8536 4564
rect 7472 4480 7524 4486
rect 7472 4422 7524 4428
rect 8024 4480 8076 4486
rect 8024 4422 8076 4428
rect 7484 4146 7512 4422
rect 8036 4214 8064 4422
rect 8214 4380 8522 4389
rect 8214 4378 8220 4380
rect 8276 4378 8300 4380
rect 8356 4378 8380 4380
rect 8436 4378 8460 4380
rect 8516 4378 8522 4380
rect 8276 4326 8278 4378
rect 8458 4326 8460 4378
rect 8214 4324 8220 4326
rect 8276 4324 8300 4326
rect 8356 4324 8380 4326
rect 8436 4324 8460 4326
rect 8516 4324 8522 4326
rect 8214 4315 8522 4324
rect 8024 4208 8076 4214
rect 8024 4150 8076 4156
rect 8680 4146 8708 6054
rect 8760 5704 8812 5710
rect 8864 5692 8892 6258
rect 8944 5840 8996 5846
rect 8944 5782 8996 5788
rect 8812 5664 8892 5692
rect 8760 5646 8812 5652
rect 7472 4140 7524 4146
rect 7472 4082 7524 4088
rect 8116 4140 8168 4146
rect 8116 4082 8168 4088
rect 8576 4140 8628 4146
rect 8576 4082 8628 4088
rect 8668 4140 8720 4146
rect 8668 4082 8720 4088
rect 7472 3936 7524 3942
rect 7472 3878 7524 3884
rect 7564 3936 7616 3942
rect 7564 3878 7616 3884
rect 7380 3732 7432 3738
rect 7380 3674 7432 3680
rect 7484 3670 7512 3878
rect 7472 3664 7524 3670
rect 7472 3606 7524 3612
rect 7576 3534 7604 3878
rect 7564 3528 7616 3534
rect 7564 3470 7616 3476
rect 7748 3528 7800 3534
rect 7748 3470 7800 3476
rect 7564 3052 7616 3058
rect 7564 2994 7616 3000
rect 7380 2984 7432 2990
rect 7380 2926 7432 2932
rect 7196 2916 7248 2922
rect 7196 2858 7248 2864
rect 7024 2746 7144 2774
rect 7024 2514 7052 2746
rect 7208 2514 7236 2858
rect 7288 2848 7340 2854
rect 7288 2790 7340 2796
rect 7012 2508 7064 2514
rect 7012 2450 7064 2456
rect 7196 2508 7248 2514
rect 7196 2450 7248 2456
rect 6736 2372 6788 2378
rect 6736 2314 6788 2320
rect 6828 2304 6880 2310
rect 6828 2246 6880 2252
rect 6736 1896 6788 1902
rect 6736 1838 6788 1844
rect 6748 1358 6776 1838
rect 6840 1562 6868 2246
rect 7300 1970 7328 2790
rect 7392 2428 7420 2926
rect 7472 2440 7524 2446
rect 7392 2400 7472 2428
rect 7472 2382 7524 2388
rect 7288 1964 7340 1970
rect 7288 1906 7340 1912
rect 7484 1902 7512 2382
rect 7576 1970 7604 2994
rect 7760 2106 7788 3470
rect 8128 3194 8156 4082
rect 8300 4004 8352 4010
rect 8300 3946 8352 3952
rect 8312 3534 8340 3946
rect 8300 3528 8352 3534
rect 8300 3470 8352 3476
rect 8214 3292 8522 3301
rect 8214 3290 8220 3292
rect 8276 3290 8300 3292
rect 8356 3290 8380 3292
rect 8436 3290 8460 3292
rect 8516 3290 8522 3292
rect 8276 3238 8278 3290
rect 8458 3238 8460 3290
rect 8214 3236 8220 3238
rect 8276 3236 8300 3238
rect 8356 3236 8380 3238
rect 8436 3236 8460 3238
rect 8516 3236 8522 3238
rect 8214 3227 8522 3236
rect 8116 3188 8168 3194
rect 8116 3130 8168 3136
rect 8588 2650 8616 4082
rect 8772 4010 8800 5646
rect 8956 5370 8984 5782
rect 9048 5710 9076 7278
rect 9324 6662 9352 8366
rect 9416 6934 9444 10406
rect 9508 10130 9536 10474
rect 9496 10124 9548 10130
rect 9496 10066 9548 10072
rect 9680 10124 9732 10130
rect 9680 10066 9732 10072
rect 9588 9376 9640 9382
rect 9588 9318 9640 9324
rect 9600 9042 9628 9318
rect 9588 9036 9640 9042
rect 9588 8978 9640 8984
rect 9692 8820 9720 10066
rect 9876 9654 9904 10610
rect 9864 9648 9916 9654
rect 9864 9590 9916 9596
rect 9692 8792 9812 8820
rect 9680 8492 9732 8498
rect 9680 8434 9732 8440
rect 9692 8022 9720 8434
rect 9784 8430 9812 8792
rect 9772 8424 9824 8430
rect 9772 8366 9824 8372
rect 9680 8016 9732 8022
rect 9680 7958 9732 7964
rect 9784 7954 9812 8366
rect 9772 7948 9824 7954
rect 9772 7890 9824 7896
rect 9588 7472 9640 7478
rect 9588 7414 9640 7420
rect 9496 7200 9548 7206
rect 9496 7142 9548 7148
rect 9404 6928 9456 6934
rect 9404 6870 9456 6876
rect 9312 6656 9364 6662
rect 9312 6598 9364 6604
rect 9324 6390 9352 6598
rect 9220 6384 9272 6390
rect 9220 6326 9272 6332
rect 9312 6384 9364 6390
rect 9312 6326 9364 6332
rect 9036 5704 9088 5710
rect 9036 5646 9088 5652
rect 8944 5364 8996 5370
rect 8944 5306 8996 5312
rect 9128 5296 9180 5302
rect 9128 5238 9180 5244
rect 9140 4826 9168 5238
rect 9128 4820 9180 4826
rect 9128 4762 9180 4768
rect 9128 4140 9180 4146
rect 9128 4082 9180 4088
rect 8760 4004 8812 4010
rect 8760 3946 8812 3952
rect 9140 3942 9168 4082
rect 9232 4078 9260 6326
rect 9324 4622 9352 6326
rect 9416 6202 9444 6870
rect 9508 6866 9536 7142
rect 9600 6866 9628 7414
rect 9784 7002 9812 7890
rect 10152 7818 10180 12310
rect 10324 11756 10376 11762
rect 10324 11698 10376 11704
rect 10336 10810 10364 11698
rect 10428 11218 10456 13330
rect 10520 12986 10548 13670
rect 10796 12986 10824 14282
rect 11060 14272 11112 14278
rect 11060 14214 11112 14220
rect 11244 14272 11296 14278
rect 11244 14214 11296 14220
rect 11980 14272 12032 14278
rect 11980 14214 12032 14220
rect 11072 13938 11100 14214
rect 11060 13932 11112 13938
rect 11060 13874 11112 13880
rect 10876 13728 10928 13734
rect 10876 13670 10928 13676
rect 10508 12980 10560 12986
rect 10508 12922 10560 12928
rect 10784 12980 10836 12986
rect 10784 12922 10836 12928
rect 10888 12850 10916 13670
rect 11072 12918 11100 13874
rect 11256 13870 11284 14214
rect 11992 13870 12020 14214
rect 12084 13870 12112 14962
rect 12716 14884 12768 14890
rect 12716 14826 12768 14832
rect 12624 14816 12676 14822
rect 12624 14758 12676 14764
rect 12214 14716 12522 14725
rect 12214 14714 12220 14716
rect 12276 14714 12300 14716
rect 12356 14714 12380 14716
rect 12436 14714 12460 14716
rect 12516 14714 12522 14716
rect 12276 14662 12278 14714
rect 12458 14662 12460 14714
rect 12214 14660 12220 14662
rect 12276 14660 12300 14662
rect 12356 14660 12380 14662
rect 12436 14660 12460 14662
rect 12516 14660 12522 14662
rect 12214 14651 12522 14660
rect 12636 14618 12664 14758
rect 12624 14612 12676 14618
rect 12624 14554 12676 14560
rect 12728 14414 12756 14826
rect 12716 14408 12768 14414
rect 12716 14350 12768 14356
rect 12808 14408 12860 14414
rect 12808 14350 12860 14356
rect 12900 14408 12952 14414
rect 12900 14350 12952 14356
rect 12624 14340 12676 14346
rect 12624 14282 12676 14288
rect 12636 13870 12664 14282
rect 11152 13864 11204 13870
rect 11152 13806 11204 13812
rect 11244 13864 11296 13870
rect 11244 13806 11296 13812
rect 11980 13864 12032 13870
rect 11980 13806 12032 13812
rect 12072 13864 12124 13870
rect 12072 13806 12124 13812
rect 12624 13864 12676 13870
rect 12624 13806 12676 13812
rect 11164 12986 11192 13806
rect 11152 12980 11204 12986
rect 11152 12922 11204 12928
rect 11060 12912 11112 12918
rect 11060 12854 11112 12860
rect 10876 12844 10928 12850
rect 10876 12786 10928 12792
rect 10888 12442 10916 12786
rect 11256 12714 11284 13806
rect 12084 13530 12112 13806
rect 12214 13628 12522 13637
rect 12214 13626 12220 13628
rect 12276 13626 12300 13628
rect 12356 13626 12380 13628
rect 12436 13626 12460 13628
rect 12516 13626 12522 13628
rect 12276 13574 12278 13626
rect 12458 13574 12460 13626
rect 12214 13572 12220 13574
rect 12276 13572 12300 13574
rect 12356 13572 12380 13574
rect 12436 13572 12460 13574
rect 12516 13572 12522 13574
rect 12214 13563 12522 13572
rect 12072 13524 12124 13530
rect 12072 13466 12124 13472
rect 12820 13394 12848 14350
rect 12912 13938 12940 14350
rect 13096 14346 13124 15370
rect 13188 15094 13216 15370
rect 13176 15088 13228 15094
rect 13176 15030 13228 15036
rect 13188 14346 13216 15030
rect 13648 14890 13676 15438
rect 13728 15020 13780 15026
rect 13728 14962 13780 14968
rect 13636 14884 13688 14890
rect 13636 14826 13688 14832
rect 13740 14618 13768 14962
rect 15120 14958 15148 16050
rect 15108 14952 15160 14958
rect 15108 14894 15160 14900
rect 13728 14612 13780 14618
rect 13728 14554 13780 14560
rect 14464 14476 14516 14482
rect 14464 14418 14516 14424
rect 13268 14408 13320 14414
rect 13268 14350 13320 14356
rect 14188 14408 14240 14414
rect 14188 14350 14240 14356
rect 13084 14340 13136 14346
rect 13084 14282 13136 14288
rect 13176 14340 13228 14346
rect 13176 14282 13228 14288
rect 12900 13932 12952 13938
rect 12900 13874 12952 13880
rect 13280 13394 13308 14350
rect 14096 13932 14148 13938
rect 14096 13874 14148 13880
rect 13360 13728 13412 13734
rect 13360 13670 13412 13676
rect 12808 13388 12860 13394
rect 12808 13330 12860 13336
rect 13268 13388 13320 13394
rect 13268 13330 13320 13336
rect 13372 13326 13400 13670
rect 14108 13394 14136 13874
rect 14200 13530 14228 14350
rect 14372 14272 14424 14278
rect 14372 14214 14424 14220
rect 14384 14006 14412 14214
rect 14372 14000 14424 14006
rect 14372 13942 14424 13948
rect 14188 13524 14240 13530
rect 14188 13466 14240 13472
rect 14476 13394 14504 14418
rect 15120 13870 15148 14894
rect 15108 13864 15160 13870
rect 15108 13806 15160 13812
rect 15396 13802 15424 16458
rect 15580 16182 15608 17614
rect 15936 17604 15988 17610
rect 15936 17546 15988 17552
rect 15752 16584 15804 16590
rect 15752 16526 15804 16532
rect 15568 16176 15620 16182
rect 15568 16118 15620 16124
rect 15764 14618 15792 16526
rect 15752 14612 15804 14618
rect 15752 14554 15804 14560
rect 15752 14408 15804 14414
rect 15752 14350 15804 14356
rect 15844 14408 15896 14414
rect 15844 14350 15896 14356
rect 15476 13932 15528 13938
rect 15476 13874 15528 13880
rect 15384 13796 15436 13802
rect 15384 13738 15436 13744
rect 14096 13388 14148 13394
rect 14096 13330 14148 13336
rect 14464 13388 14516 13394
rect 14464 13330 14516 13336
rect 13360 13320 13412 13326
rect 13360 13262 13412 13268
rect 13634 12880 13690 12889
rect 13634 12815 13690 12824
rect 11244 12708 11296 12714
rect 11244 12650 11296 12656
rect 12214 12540 12522 12549
rect 12214 12538 12220 12540
rect 12276 12538 12300 12540
rect 12356 12538 12380 12540
rect 12436 12538 12460 12540
rect 12516 12538 12522 12540
rect 12276 12486 12278 12538
rect 12458 12486 12460 12538
rect 12214 12484 12220 12486
rect 12276 12484 12300 12486
rect 12356 12484 12380 12486
rect 12436 12484 12460 12486
rect 12516 12484 12522 12486
rect 12214 12475 12522 12484
rect 10876 12436 10928 12442
rect 10876 12378 10928 12384
rect 11796 12300 11848 12306
rect 11796 12242 11848 12248
rect 11244 12232 11296 12238
rect 10690 12200 10746 12209
rect 11244 12174 11296 12180
rect 11520 12232 11572 12238
rect 11520 12174 11572 12180
rect 10690 12135 10746 12144
rect 10704 11898 10732 12135
rect 11256 11898 11284 12174
rect 10692 11892 10744 11898
rect 10692 11834 10744 11840
rect 11244 11892 11296 11898
rect 11244 11834 11296 11840
rect 11428 11620 11480 11626
rect 11428 11562 11480 11568
rect 11440 11354 11468 11562
rect 11428 11348 11480 11354
rect 11428 11290 11480 11296
rect 10416 11212 10468 11218
rect 10416 11154 10468 11160
rect 10324 10804 10376 10810
rect 10324 10746 10376 10752
rect 10324 10600 10376 10606
rect 10324 10542 10376 10548
rect 10336 10198 10364 10542
rect 10324 10192 10376 10198
rect 10324 10134 10376 10140
rect 10428 10130 10456 11154
rect 11060 11144 11112 11150
rect 11060 11086 11112 11092
rect 10784 10668 10836 10674
rect 10784 10610 10836 10616
rect 10796 10470 10824 10610
rect 10784 10464 10836 10470
rect 10784 10406 10836 10412
rect 10416 10124 10468 10130
rect 10416 10066 10468 10072
rect 10692 9988 10744 9994
rect 10692 9930 10744 9936
rect 10704 9722 10732 9930
rect 10692 9716 10744 9722
rect 10692 9658 10744 9664
rect 10784 9648 10836 9654
rect 10784 9590 10836 9596
rect 10416 9580 10468 9586
rect 10416 9522 10468 9528
rect 10692 9580 10744 9586
rect 10692 9522 10744 9528
rect 10428 8634 10456 9522
rect 10600 8900 10652 8906
rect 10600 8842 10652 8848
rect 10612 8634 10640 8842
rect 10416 8628 10468 8634
rect 10416 8570 10468 8576
rect 10600 8628 10652 8634
rect 10600 8570 10652 8576
rect 10600 8424 10652 8430
rect 10600 8366 10652 8372
rect 10140 7812 10192 7818
rect 10140 7754 10192 7760
rect 10152 7410 10180 7754
rect 10140 7404 10192 7410
rect 10140 7346 10192 7352
rect 9956 7200 10008 7206
rect 9956 7142 10008 7148
rect 9772 6996 9824 7002
rect 9772 6938 9824 6944
rect 9496 6860 9548 6866
rect 9496 6802 9548 6808
rect 9588 6860 9640 6866
rect 9588 6802 9640 6808
rect 9416 6186 9536 6202
rect 9784 6186 9812 6938
rect 9968 6798 9996 7142
rect 9956 6792 10008 6798
rect 9956 6734 10008 6740
rect 9968 6322 9996 6734
rect 10508 6452 10560 6458
rect 10508 6394 10560 6400
rect 9864 6316 9916 6322
rect 9864 6258 9916 6264
rect 9956 6316 10008 6322
rect 9956 6258 10008 6264
rect 9404 6180 9536 6186
rect 9456 6174 9536 6180
rect 9404 6122 9456 6128
rect 9508 5574 9536 6174
rect 9772 6180 9824 6186
rect 9772 6122 9824 6128
rect 9588 6112 9640 6118
rect 9588 6054 9640 6060
rect 9496 5568 9548 5574
rect 9496 5510 9548 5516
rect 9600 5302 9628 6054
rect 9876 5370 9904 6258
rect 9864 5364 9916 5370
rect 9864 5306 9916 5312
rect 9588 5296 9640 5302
rect 9588 5238 9640 5244
rect 9968 4622 9996 6258
rect 10324 6248 10376 6254
rect 10324 6190 10376 6196
rect 10048 6112 10100 6118
rect 10048 6054 10100 6060
rect 10060 5642 10088 6054
rect 10048 5636 10100 5642
rect 10048 5578 10100 5584
rect 10336 5234 10364 6190
rect 10324 5228 10376 5234
rect 10324 5170 10376 5176
rect 10520 4758 10548 6394
rect 10508 4752 10560 4758
rect 10508 4694 10560 4700
rect 9312 4616 9364 4622
rect 9312 4558 9364 4564
rect 9956 4616 10008 4622
rect 9956 4558 10008 4564
rect 10520 4282 10548 4694
rect 10508 4276 10560 4282
rect 10508 4218 10560 4224
rect 9220 4072 9272 4078
rect 9220 4014 9272 4020
rect 9128 3936 9180 3942
rect 9128 3878 9180 3884
rect 8852 3732 8904 3738
rect 8852 3674 8904 3680
rect 8576 2644 8628 2650
rect 8576 2586 8628 2592
rect 8116 2304 8168 2310
rect 8116 2246 8168 2252
rect 7748 2100 7800 2106
rect 7748 2042 7800 2048
rect 7564 1964 7616 1970
rect 7564 1906 7616 1912
rect 7380 1896 7432 1902
rect 7380 1838 7432 1844
rect 7472 1896 7524 1902
rect 7472 1838 7524 1844
rect 6828 1556 6880 1562
rect 6828 1498 6880 1504
rect 7392 1426 7420 1838
rect 8128 1426 8156 2246
rect 8214 2204 8522 2213
rect 8214 2202 8220 2204
rect 8276 2202 8300 2204
rect 8356 2202 8380 2204
rect 8436 2202 8460 2204
rect 8516 2202 8522 2204
rect 8276 2150 8278 2202
rect 8458 2150 8460 2202
rect 8214 2148 8220 2150
rect 8276 2148 8300 2150
rect 8356 2148 8380 2150
rect 8436 2148 8460 2150
rect 8516 2148 8522 2150
rect 8214 2139 8522 2148
rect 8668 1964 8720 1970
rect 8668 1906 8720 1912
rect 8392 1896 8444 1902
rect 8392 1838 8444 1844
rect 8404 1562 8432 1838
rect 8392 1556 8444 1562
rect 8392 1498 8444 1504
rect 8680 1494 8708 1906
rect 8864 1766 8892 3674
rect 9036 3596 9088 3602
rect 9036 3538 9088 3544
rect 9048 3058 9076 3538
rect 9036 3052 9088 3058
rect 9036 2994 9088 3000
rect 9140 2446 9168 3878
rect 9232 3466 9260 4014
rect 9772 3936 9824 3942
rect 9772 3878 9824 3884
rect 9784 3466 9812 3878
rect 10520 3738 10548 4218
rect 10612 4146 10640 8366
rect 10704 8090 10732 9522
rect 10796 8498 10824 9590
rect 11072 9450 11100 11086
rect 11244 11008 11296 11014
rect 11244 10950 11296 10956
rect 11152 10464 11204 10470
rect 11152 10406 11204 10412
rect 11060 9444 11112 9450
rect 11060 9386 11112 9392
rect 11164 9178 11192 10406
rect 11256 10130 11284 10950
rect 11440 10810 11468 11290
rect 11532 10810 11560 12174
rect 11704 12096 11756 12102
rect 11704 12038 11756 12044
rect 11716 11354 11744 12038
rect 11808 11898 11836 12242
rect 13648 12238 13676 12815
rect 13636 12232 13688 12238
rect 13636 12174 13688 12180
rect 11796 11892 11848 11898
rect 11796 11834 11848 11840
rect 12808 11620 12860 11626
rect 12808 11562 12860 11568
rect 13360 11620 13412 11626
rect 13360 11562 13412 11568
rect 12214 11452 12522 11461
rect 12214 11450 12220 11452
rect 12276 11450 12300 11452
rect 12356 11450 12380 11452
rect 12436 11450 12460 11452
rect 12516 11450 12522 11452
rect 12276 11398 12278 11450
rect 12458 11398 12460 11450
rect 12214 11396 12220 11398
rect 12276 11396 12300 11398
rect 12356 11396 12380 11398
rect 12436 11396 12460 11398
rect 12516 11396 12522 11398
rect 12214 11387 12522 11396
rect 11704 11348 11756 11354
rect 11704 11290 11756 11296
rect 12164 11348 12216 11354
rect 12164 11290 12216 11296
rect 11428 10804 11480 10810
rect 11428 10746 11480 10752
rect 11520 10804 11572 10810
rect 11520 10746 11572 10752
rect 11336 10668 11388 10674
rect 11336 10610 11388 10616
rect 11244 10124 11296 10130
rect 11244 10066 11296 10072
rect 11256 9586 11284 10066
rect 11244 9580 11296 9586
rect 11244 9522 11296 9528
rect 11152 9172 11204 9178
rect 11152 9114 11204 9120
rect 10784 8492 10836 8498
rect 10784 8434 10836 8440
rect 10692 8084 10744 8090
rect 10692 8026 10744 8032
rect 11164 7954 11192 9114
rect 11256 8498 11284 9522
rect 11244 8492 11296 8498
rect 11244 8434 11296 8440
rect 11152 7948 11204 7954
rect 11152 7890 11204 7896
rect 11060 7540 11112 7546
rect 11060 7482 11112 7488
rect 10968 6860 11020 6866
rect 10968 6802 11020 6808
rect 10980 5234 11008 6802
rect 11072 6662 11100 7482
rect 11060 6656 11112 6662
rect 11060 6598 11112 6604
rect 10968 5228 11020 5234
rect 10968 5170 11020 5176
rect 10980 4282 11008 5170
rect 11152 4752 11204 4758
rect 11152 4694 11204 4700
rect 10968 4276 11020 4282
rect 10968 4218 11020 4224
rect 10600 4140 10652 4146
rect 10600 4082 10652 4088
rect 10600 3936 10652 3942
rect 10600 3878 10652 3884
rect 10508 3732 10560 3738
rect 10508 3674 10560 3680
rect 9864 3596 9916 3602
rect 9864 3538 9916 3544
rect 9220 3460 9272 3466
rect 9220 3402 9272 3408
rect 9772 3460 9824 3466
rect 9772 3402 9824 3408
rect 9232 2836 9260 3402
rect 9312 3392 9364 3398
rect 9312 3334 9364 3340
rect 9324 3126 9352 3334
rect 9496 3188 9548 3194
rect 9496 3130 9548 3136
rect 9312 3120 9364 3126
rect 9312 3062 9364 3068
rect 9404 2984 9456 2990
rect 9508 2938 9536 3130
rect 9456 2932 9536 2938
rect 9404 2926 9536 2932
rect 9416 2910 9536 2926
rect 9312 2848 9364 2854
rect 9232 2808 9312 2836
rect 9128 2440 9180 2446
rect 9128 2382 9180 2388
rect 9232 1902 9260 2808
rect 9312 2790 9364 2796
rect 9508 2106 9536 2910
rect 9876 2514 9904 3538
rect 10612 3534 10640 3878
rect 10980 3602 11008 4218
rect 11164 4146 11192 4694
rect 11152 4140 11204 4146
rect 11152 4082 11204 4088
rect 11348 4010 11376 10610
rect 12176 10538 12204 11290
rect 12624 11076 12676 11082
rect 12624 11018 12676 11024
rect 12348 10736 12400 10742
rect 12348 10678 12400 10684
rect 12164 10532 12216 10538
rect 12164 10474 12216 10480
rect 12360 10470 12388 10678
rect 12348 10464 12400 10470
rect 12348 10406 12400 10412
rect 12214 10364 12522 10373
rect 12214 10362 12220 10364
rect 12276 10362 12300 10364
rect 12356 10362 12380 10364
rect 12436 10362 12460 10364
rect 12516 10362 12522 10364
rect 12276 10310 12278 10362
rect 12458 10310 12460 10362
rect 12214 10308 12220 10310
rect 12276 10308 12300 10310
rect 12356 10308 12380 10310
rect 12436 10308 12460 10310
rect 12516 10308 12522 10310
rect 12214 10299 12522 10308
rect 12636 10266 12664 11018
rect 12716 11008 12768 11014
rect 12716 10950 12768 10956
rect 12728 10810 12756 10950
rect 12716 10804 12768 10810
rect 12716 10746 12768 10752
rect 12716 10668 12768 10674
rect 12820 10656 12848 11562
rect 13372 10810 13400 11562
rect 13648 11150 13676 12174
rect 14108 11914 14136 13330
rect 15016 13252 15068 13258
rect 15016 13194 15068 13200
rect 15028 12986 15056 13194
rect 15488 12986 15516 13874
rect 15764 13530 15792 14350
rect 15856 13870 15884 14350
rect 15844 13864 15896 13870
rect 15844 13806 15896 13812
rect 15752 13524 15804 13530
rect 15752 13466 15804 13472
rect 15016 12980 15068 12986
rect 15016 12922 15068 12928
rect 15476 12980 15528 12986
rect 15476 12922 15528 12928
rect 15016 12844 15068 12850
rect 15016 12786 15068 12792
rect 14832 12776 14884 12782
rect 14832 12718 14884 12724
rect 14844 12238 14872 12718
rect 15028 12238 15056 12786
rect 15568 12300 15620 12306
rect 15568 12242 15620 12248
rect 14832 12232 14884 12238
rect 14832 12174 14884 12180
rect 15016 12232 15068 12238
rect 15016 12174 15068 12180
rect 14016 11898 14136 11914
rect 13820 11892 13872 11898
rect 13820 11834 13872 11840
rect 14004 11892 14136 11898
rect 14056 11886 14136 11892
rect 14280 11892 14332 11898
rect 14004 11834 14056 11840
rect 14280 11834 14332 11840
rect 13636 11144 13688 11150
rect 13636 11086 13688 11092
rect 13832 11082 13860 11834
rect 14016 11218 14044 11834
rect 14292 11354 14320 11834
rect 14844 11354 14872 12174
rect 14924 12096 14976 12102
rect 14924 12038 14976 12044
rect 14936 11830 14964 12038
rect 14924 11824 14976 11830
rect 14924 11766 14976 11772
rect 15108 11552 15160 11558
rect 15108 11494 15160 11500
rect 14280 11348 14332 11354
rect 14280 11290 14332 11296
rect 14832 11348 14884 11354
rect 14832 11290 14884 11296
rect 14004 11212 14056 11218
rect 14004 11154 14056 11160
rect 13820 11076 13872 11082
rect 13820 11018 13872 11024
rect 14740 11076 14792 11082
rect 14740 11018 14792 11024
rect 13728 11008 13780 11014
rect 13728 10950 13780 10956
rect 13740 10810 13768 10950
rect 13360 10804 13412 10810
rect 13360 10746 13412 10752
rect 13728 10804 13780 10810
rect 13728 10746 13780 10752
rect 12900 10736 12952 10742
rect 12900 10678 12952 10684
rect 12768 10628 12848 10656
rect 12716 10610 12768 10616
rect 12624 10260 12676 10266
rect 12624 10202 12676 10208
rect 12728 10062 12756 10610
rect 12912 10130 12940 10678
rect 14464 10464 14516 10470
rect 14464 10406 14516 10412
rect 12900 10124 12952 10130
rect 12900 10066 12952 10072
rect 12716 10056 12768 10062
rect 12716 9998 12768 10004
rect 11980 9988 12032 9994
rect 11980 9930 12032 9936
rect 11704 9920 11756 9926
rect 11704 9862 11756 9868
rect 11716 9654 11744 9862
rect 11992 9654 12020 9930
rect 12164 9920 12216 9926
rect 12164 9862 12216 9868
rect 11704 9648 11756 9654
rect 11704 9590 11756 9596
rect 11980 9648 12032 9654
rect 11980 9590 12032 9596
rect 11520 9376 11572 9382
rect 11520 9318 11572 9324
rect 11532 8566 11560 9318
rect 11716 8922 11744 9590
rect 12072 9580 12124 9586
rect 12072 9522 12124 9528
rect 11716 8894 11836 8922
rect 11704 8832 11756 8838
rect 11704 8774 11756 8780
rect 11520 8560 11572 8566
rect 11520 8502 11572 8508
rect 11716 8430 11744 8774
rect 11704 8424 11756 8430
rect 11704 8366 11756 8372
rect 11808 7818 11836 8894
rect 11888 8900 11940 8906
rect 11888 8842 11940 8848
rect 11900 8634 11928 8842
rect 11888 8628 11940 8634
rect 11888 8570 11940 8576
rect 11888 8492 11940 8498
rect 11888 8434 11940 8440
rect 11980 8492 12032 8498
rect 11980 8434 12032 8440
rect 11900 8090 11928 8434
rect 11888 8084 11940 8090
rect 11888 8026 11940 8032
rect 11796 7812 11848 7818
rect 11796 7754 11848 7760
rect 11992 7410 12020 8434
rect 12084 7886 12112 9522
rect 12176 9382 12204 9862
rect 12164 9376 12216 9382
rect 12164 9318 12216 9324
rect 12214 9276 12522 9285
rect 12214 9274 12220 9276
rect 12276 9274 12300 9276
rect 12356 9274 12380 9276
rect 12436 9274 12460 9276
rect 12516 9274 12522 9276
rect 12276 9222 12278 9274
rect 12458 9222 12460 9274
rect 12214 9220 12220 9222
rect 12276 9220 12300 9222
rect 12356 9220 12380 9222
rect 12436 9220 12460 9222
rect 12516 9220 12522 9222
rect 12214 9211 12522 9220
rect 12440 8832 12492 8838
rect 12440 8774 12492 8780
rect 12452 8634 12480 8774
rect 12440 8628 12492 8634
rect 12440 8570 12492 8576
rect 12214 8188 12522 8197
rect 12214 8186 12220 8188
rect 12276 8186 12300 8188
rect 12356 8186 12380 8188
rect 12436 8186 12460 8188
rect 12516 8186 12522 8188
rect 12276 8134 12278 8186
rect 12458 8134 12460 8186
rect 12214 8132 12220 8134
rect 12276 8132 12300 8134
rect 12356 8132 12380 8134
rect 12436 8132 12460 8134
rect 12516 8132 12522 8134
rect 12214 8123 12522 8132
rect 12256 8084 12308 8090
rect 12256 8026 12308 8032
rect 12072 7880 12124 7886
rect 12072 7822 12124 7828
rect 12268 7410 12296 8026
rect 11796 7404 11848 7410
rect 11796 7346 11848 7352
rect 11980 7404 12032 7410
rect 11980 7346 12032 7352
rect 12256 7404 12308 7410
rect 12256 7346 12308 7352
rect 11612 7200 11664 7206
rect 11612 7142 11664 7148
rect 11624 7002 11652 7142
rect 11612 6996 11664 7002
rect 11612 6938 11664 6944
rect 11808 6458 11836 7346
rect 11980 7200 12032 7206
rect 11980 7142 12032 7148
rect 11992 6730 12020 7142
rect 12214 7100 12522 7109
rect 12214 7098 12220 7100
rect 12276 7098 12300 7100
rect 12356 7098 12380 7100
rect 12436 7098 12460 7100
rect 12516 7098 12522 7100
rect 12276 7046 12278 7098
rect 12458 7046 12460 7098
rect 12214 7044 12220 7046
rect 12276 7044 12300 7046
rect 12356 7044 12380 7046
rect 12436 7044 12460 7046
rect 12516 7044 12522 7046
rect 12214 7035 12522 7044
rect 12728 6914 12756 9998
rect 13084 9920 13136 9926
rect 13084 9862 13136 9868
rect 12900 7744 12952 7750
rect 12900 7686 12952 7692
rect 12912 7478 12940 7686
rect 12900 7472 12952 7478
rect 12900 7414 12952 7420
rect 12636 6886 12756 6914
rect 12440 6860 12492 6866
rect 12440 6802 12492 6808
rect 12452 6746 12480 6802
rect 12636 6798 12664 6886
rect 11980 6724 12032 6730
rect 11980 6666 12032 6672
rect 12084 6718 12480 6746
rect 12624 6792 12676 6798
rect 12624 6734 12676 6740
rect 11796 6452 11848 6458
rect 11796 6394 11848 6400
rect 11428 6316 11480 6322
rect 11428 6258 11480 6264
rect 11440 5914 11468 6258
rect 12084 5914 12112 6718
rect 12256 6656 12308 6662
rect 12256 6598 12308 6604
rect 12268 6458 12296 6598
rect 12256 6452 12308 6458
rect 12256 6394 12308 6400
rect 12636 6390 12664 6734
rect 12624 6384 12676 6390
rect 12624 6326 12676 6332
rect 12214 6012 12522 6021
rect 12214 6010 12220 6012
rect 12276 6010 12300 6012
rect 12356 6010 12380 6012
rect 12436 6010 12460 6012
rect 12516 6010 12522 6012
rect 12276 5958 12278 6010
rect 12458 5958 12460 6010
rect 12214 5956 12220 5958
rect 12276 5956 12300 5958
rect 12356 5956 12380 5958
rect 12436 5956 12460 5958
rect 12516 5956 12522 5958
rect 12214 5947 12522 5956
rect 11428 5908 11480 5914
rect 11428 5850 11480 5856
rect 12072 5908 12124 5914
rect 12072 5850 12124 5856
rect 11440 5710 11468 5850
rect 11428 5704 11480 5710
rect 11426 5672 11428 5681
rect 11480 5672 11482 5681
rect 11426 5607 11482 5616
rect 11980 5636 12032 5642
rect 11980 5578 12032 5584
rect 11520 5568 11572 5574
rect 11520 5510 11572 5516
rect 11428 4616 11480 4622
rect 11428 4558 11480 4564
rect 11336 4004 11388 4010
rect 11336 3946 11388 3952
rect 11152 3936 11204 3942
rect 11152 3878 11204 3884
rect 10968 3596 11020 3602
rect 10968 3538 11020 3544
rect 10600 3528 10652 3534
rect 10600 3470 10652 3476
rect 11164 3126 11192 3878
rect 11348 3738 11376 3946
rect 11440 3942 11468 4558
rect 11532 4486 11560 5510
rect 11888 5160 11940 5166
rect 11888 5102 11940 5108
rect 11900 4826 11928 5102
rect 11992 5030 12020 5578
rect 12072 5568 12124 5574
rect 12072 5510 12124 5516
rect 11980 5024 12032 5030
rect 11980 4966 12032 4972
rect 11888 4820 11940 4826
rect 11888 4762 11940 4768
rect 11992 4690 12020 4966
rect 11980 4684 12032 4690
rect 11980 4626 12032 4632
rect 12084 4622 12112 5510
rect 12624 5296 12676 5302
rect 12624 5238 12676 5244
rect 12214 4924 12522 4933
rect 12214 4922 12220 4924
rect 12276 4922 12300 4924
rect 12356 4922 12380 4924
rect 12436 4922 12460 4924
rect 12516 4922 12522 4924
rect 12276 4870 12278 4922
rect 12458 4870 12460 4922
rect 12214 4868 12220 4870
rect 12276 4868 12300 4870
rect 12356 4868 12380 4870
rect 12436 4868 12460 4870
rect 12516 4868 12522 4870
rect 12214 4859 12522 4868
rect 12636 4826 12664 5238
rect 12624 4820 12676 4826
rect 12624 4762 12676 4768
rect 12072 4616 12124 4622
rect 12072 4558 12124 4564
rect 12624 4548 12676 4554
rect 12624 4490 12676 4496
rect 11520 4480 11572 4486
rect 11520 4422 11572 4428
rect 11980 4072 12032 4078
rect 11980 4014 12032 4020
rect 11428 3936 11480 3942
rect 11428 3878 11480 3884
rect 11992 3738 12020 4014
rect 12214 3836 12522 3845
rect 12214 3834 12220 3836
rect 12276 3834 12300 3836
rect 12356 3834 12380 3836
rect 12436 3834 12460 3836
rect 12516 3834 12522 3836
rect 12276 3782 12278 3834
rect 12458 3782 12460 3834
rect 12214 3780 12220 3782
rect 12276 3780 12300 3782
rect 12356 3780 12380 3782
rect 12436 3780 12460 3782
rect 12516 3780 12522 3782
rect 12214 3771 12522 3780
rect 11336 3732 11388 3738
rect 11336 3674 11388 3680
rect 11980 3732 12032 3738
rect 11980 3674 12032 3680
rect 12072 3460 12124 3466
rect 12072 3402 12124 3408
rect 11152 3120 11204 3126
rect 11152 3062 11204 3068
rect 12084 2922 12112 3402
rect 12636 3058 12664 4490
rect 12992 4480 13044 4486
rect 12992 4422 13044 4428
rect 13004 4214 13032 4422
rect 12992 4208 13044 4214
rect 12992 4150 13044 4156
rect 12992 3936 13044 3942
rect 12992 3878 13044 3884
rect 13004 3534 13032 3878
rect 13096 3670 13124 9862
rect 14476 9654 14504 10406
rect 14464 9648 14516 9654
rect 14464 9590 14516 9596
rect 13176 9512 13228 9518
rect 13176 9454 13228 9460
rect 13188 9042 13216 9454
rect 13176 9036 13228 9042
rect 13176 8978 13228 8984
rect 14556 9036 14608 9042
rect 14556 8978 14608 8984
rect 13188 7342 13216 8978
rect 14568 8378 14596 8978
rect 14476 8362 14596 8378
rect 13820 8356 13872 8362
rect 13820 8298 13872 8304
rect 14464 8356 14596 8362
rect 14516 8350 14596 8356
rect 14464 8298 14516 8304
rect 13636 7744 13688 7750
rect 13636 7686 13688 7692
rect 13648 7546 13676 7686
rect 13636 7540 13688 7546
rect 13636 7482 13688 7488
rect 13176 7336 13228 7342
rect 13176 7278 13228 7284
rect 13452 7336 13504 7342
rect 13452 7278 13504 7284
rect 13188 6934 13216 7278
rect 13464 7002 13492 7278
rect 13452 6996 13504 7002
rect 13452 6938 13504 6944
rect 13176 6928 13228 6934
rect 13176 6870 13228 6876
rect 13360 6384 13412 6390
rect 13360 6326 13412 6332
rect 13268 5772 13320 5778
rect 13268 5714 13320 5720
rect 13084 3664 13136 3670
rect 13084 3606 13136 3612
rect 12992 3528 13044 3534
rect 12992 3470 13044 3476
rect 13096 3058 13124 3606
rect 13280 3602 13308 5714
rect 13372 5642 13400 6326
rect 13648 5846 13676 7482
rect 13728 6656 13780 6662
rect 13728 6598 13780 6604
rect 13740 5846 13768 6598
rect 13832 6254 13860 8298
rect 14568 8090 14596 8350
rect 14556 8084 14608 8090
rect 14556 8026 14608 8032
rect 14752 7886 14780 11018
rect 15120 10742 15148 11494
rect 15580 11286 15608 12242
rect 15568 11280 15620 11286
rect 15568 11222 15620 11228
rect 15476 11008 15528 11014
rect 15476 10950 15528 10956
rect 15108 10736 15160 10742
rect 15108 10678 15160 10684
rect 15292 10736 15344 10742
rect 15292 10678 15344 10684
rect 14924 10668 14976 10674
rect 14924 10610 14976 10616
rect 14936 10266 14964 10610
rect 14924 10260 14976 10266
rect 14924 10202 14976 10208
rect 15120 10130 15148 10678
rect 15200 10464 15252 10470
rect 15200 10406 15252 10412
rect 15108 10124 15160 10130
rect 15108 10066 15160 10072
rect 15212 9674 15240 10406
rect 15304 10198 15332 10678
rect 15488 10674 15516 10950
rect 15476 10668 15528 10674
rect 15476 10610 15528 10616
rect 15292 10192 15344 10198
rect 15292 10134 15344 10140
rect 15384 9988 15436 9994
rect 15384 9930 15436 9936
rect 15292 9920 15344 9926
rect 15292 9862 15344 9868
rect 15304 9722 15332 9862
rect 15120 9646 15240 9674
rect 15292 9716 15344 9722
rect 15292 9658 15344 9664
rect 14832 8832 14884 8838
rect 14832 8774 14884 8780
rect 14844 8430 14872 8774
rect 15016 8560 15068 8566
rect 15016 8502 15068 8508
rect 14832 8424 14884 8430
rect 14832 8366 14884 8372
rect 14188 7880 14240 7886
rect 14188 7822 14240 7828
rect 14740 7880 14792 7886
rect 14740 7822 14792 7828
rect 14200 7546 14228 7822
rect 14188 7540 14240 7546
rect 14188 7482 14240 7488
rect 14844 6798 14872 8366
rect 15028 8090 15056 8502
rect 15016 8084 15068 8090
rect 15016 8026 15068 8032
rect 15120 7478 15148 9646
rect 15304 8974 15332 9658
rect 15396 8974 15424 9930
rect 15476 9648 15528 9654
rect 15476 9590 15528 9596
rect 15488 9178 15516 9590
rect 15476 9172 15528 9178
rect 15476 9114 15528 9120
rect 15292 8968 15344 8974
rect 15292 8910 15344 8916
rect 15384 8968 15436 8974
rect 15384 8910 15436 8916
rect 15476 8832 15528 8838
rect 15476 8774 15528 8780
rect 15488 8566 15516 8774
rect 15476 8560 15528 8566
rect 15476 8502 15528 8508
rect 15200 7812 15252 7818
rect 15200 7754 15252 7760
rect 15108 7472 15160 7478
rect 15108 7414 15160 7420
rect 14924 7200 14976 7206
rect 14924 7142 14976 7148
rect 14832 6792 14884 6798
rect 14832 6734 14884 6740
rect 14936 6662 14964 7142
rect 14924 6656 14976 6662
rect 14924 6598 14976 6604
rect 13912 6316 13964 6322
rect 13912 6258 13964 6264
rect 13820 6248 13872 6254
rect 13820 6190 13872 6196
rect 13636 5840 13688 5846
rect 13636 5782 13688 5788
rect 13728 5840 13780 5846
rect 13728 5782 13780 5788
rect 13360 5636 13412 5642
rect 13360 5578 13412 5584
rect 13372 5302 13400 5578
rect 13360 5296 13412 5302
rect 13360 5238 13412 5244
rect 13648 4690 13676 5782
rect 13832 5778 13860 6190
rect 13820 5772 13872 5778
rect 13820 5714 13872 5720
rect 13728 5228 13780 5234
rect 13728 5170 13780 5176
rect 13636 4684 13688 4690
rect 13636 4626 13688 4632
rect 13740 4622 13768 5170
rect 13820 5024 13872 5030
rect 13820 4966 13872 4972
rect 13832 4826 13860 4966
rect 13820 4820 13872 4826
rect 13820 4762 13872 4768
rect 13728 4616 13780 4622
rect 13728 4558 13780 4564
rect 13268 3596 13320 3602
rect 13268 3538 13320 3544
rect 12624 3052 12676 3058
rect 12624 2994 12676 3000
rect 12900 3052 12952 3058
rect 12900 2994 12952 3000
rect 13084 3052 13136 3058
rect 13820 3052 13872 3058
rect 13084 2994 13136 3000
rect 13740 3012 13820 3040
rect 12072 2916 12124 2922
rect 12072 2858 12124 2864
rect 11244 2848 11296 2854
rect 11244 2790 11296 2796
rect 9864 2508 9916 2514
rect 9864 2450 9916 2456
rect 10876 2508 10928 2514
rect 10876 2450 10928 2456
rect 9496 2100 9548 2106
rect 9496 2042 9548 2048
rect 10888 2038 10916 2450
rect 11152 2372 11204 2378
rect 11152 2314 11204 2320
rect 10876 2032 10928 2038
rect 10876 1974 10928 1980
rect 9220 1896 9272 1902
rect 9220 1838 9272 1844
rect 10968 1896 11020 1902
rect 10968 1838 11020 1844
rect 8852 1760 8904 1766
rect 8852 1702 8904 1708
rect 8668 1488 8720 1494
rect 8668 1430 8720 1436
rect 7380 1420 7432 1426
rect 7380 1362 7432 1368
rect 8116 1420 8168 1426
rect 8116 1362 8168 1368
rect 9232 1358 9260 1838
rect 10980 1562 11008 1838
rect 11164 1562 11192 2314
rect 10968 1556 11020 1562
rect 10968 1498 11020 1504
rect 11152 1556 11204 1562
rect 11152 1498 11204 1504
rect 11256 1358 11284 2790
rect 12084 1970 12112 2858
rect 12214 2748 12522 2757
rect 12214 2746 12220 2748
rect 12276 2746 12300 2748
rect 12356 2746 12380 2748
rect 12436 2746 12460 2748
rect 12516 2746 12522 2748
rect 12276 2694 12278 2746
rect 12458 2694 12460 2746
rect 12214 2692 12220 2694
rect 12276 2692 12300 2694
rect 12356 2692 12380 2694
rect 12436 2692 12460 2694
rect 12516 2692 12522 2694
rect 12214 2683 12522 2692
rect 12636 2650 12664 2994
rect 12808 2848 12860 2854
rect 12808 2790 12860 2796
rect 12624 2644 12676 2650
rect 12624 2586 12676 2592
rect 12820 2378 12848 2790
rect 12808 2372 12860 2378
rect 12808 2314 12860 2320
rect 12164 2304 12216 2310
rect 12164 2246 12216 2252
rect 12176 2106 12204 2246
rect 12164 2100 12216 2106
rect 12164 2042 12216 2048
rect 12072 1964 12124 1970
rect 12072 1906 12124 1912
rect 12176 1816 12204 2042
rect 12912 1970 12940 2994
rect 13740 2650 13768 3012
rect 13820 2994 13872 3000
rect 13728 2644 13780 2650
rect 13728 2586 13780 2592
rect 13740 2446 13768 2586
rect 13924 2514 13952 6258
rect 14464 6248 14516 6254
rect 14464 6190 14516 6196
rect 14476 5642 14504 6190
rect 14464 5636 14516 5642
rect 14464 5578 14516 5584
rect 14188 5092 14240 5098
rect 14188 5034 14240 5040
rect 14200 4146 14228 5034
rect 14476 4690 14504 5578
rect 14936 5370 14964 6598
rect 15108 6248 15160 6254
rect 15108 6190 15160 6196
rect 15120 5914 15148 6190
rect 15108 5908 15160 5914
rect 15108 5850 15160 5856
rect 14924 5364 14976 5370
rect 14924 5306 14976 5312
rect 15108 5228 15160 5234
rect 15108 5170 15160 5176
rect 14924 5160 14976 5166
rect 14924 5102 14976 5108
rect 14556 5024 14608 5030
rect 14556 4966 14608 4972
rect 14464 4684 14516 4690
rect 14464 4626 14516 4632
rect 14372 4548 14424 4554
rect 14372 4490 14424 4496
rect 14188 4140 14240 4146
rect 14188 4082 14240 4088
rect 14384 4010 14412 4490
rect 14476 4282 14504 4626
rect 14568 4554 14596 4966
rect 14556 4548 14608 4554
rect 14556 4490 14608 4496
rect 14464 4276 14516 4282
rect 14464 4218 14516 4224
rect 14476 4146 14504 4218
rect 14464 4140 14516 4146
rect 14464 4082 14516 4088
rect 14372 4004 14424 4010
rect 14372 3946 14424 3952
rect 14556 3528 14608 3534
rect 14556 3470 14608 3476
rect 14188 3392 14240 3398
rect 14188 3334 14240 3340
rect 14200 3194 14228 3334
rect 14188 3188 14240 3194
rect 14188 3130 14240 3136
rect 14200 2650 14228 3130
rect 14280 3052 14332 3058
rect 14280 2994 14332 3000
rect 14188 2644 14240 2650
rect 14188 2586 14240 2592
rect 14292 2514 14320 2994
rect 14372 2848 14424 2854
rect 14372 2790 14424 2796
rect 13912 2508 13964 2514
rect 13912 2450 13964 2456
rect 14280 2508 14332 2514
rect 14280 2450 14332 2456
rect 13084 2440 13136 2446
rect 13084 2382 13136 2388
rect 13728 2440 13780 2446
rect 13728 2382 13780 2388
rect 13096 1970 13124 2382
rect 14384 2038 14412 2790
rect 14372 2032 14424 2038
rect 14372 1974 14424 1980
rect 12900 1964 12952 1970
rect 12900 1906 12952 1912
rect 13084 1964 13136 1970
rect 13084 1906 13136 1912
rect 12084 1788 12204 1816
rect 11796 1760 11848 1766
rect 11796 1702 11848 1708
rect 11808 1358 11836 1702
rect 12084 1494 12112 1788
rect 13544 1760 13596 1766
rect 13544 1702 13596 1708
rect 12214 1660 12522 1669
rect 12214 1658 12220 1660
rect 12276 1658 12300 1660
rect 12356 1658 12380 1660
rect 12436 1658 12460 1660
rect 12516 1658 12522 1660
rect 12276 1606 12278 1658
rect 12458 1606 12460 1658
rect 12214 1604 12220 1606
rect 12276 1604 12300 1606
rect 12356 1604 12380 1606
rect 12436 1604 12460 1606
rect 12516 1604 12522 1606
rect 12214 1595 12522 1604
rect 12072 1488 12124 1494
rect 12072 1430 12124 1436
rect 13556 1358 13584 1702
rect 6736 1352 6788 1358
rect 6736 1294 6788 1300
rect 9220 1352 9272 1358
rect 9220 1294 9272 1300
rect 11244 1352 11296 1358
rect 11244 1294 11296 1300
rect 11796 1352 11848 1358
rect 11796 1294 11848 1300
rect 13544 1352 13596 1358
rect 13544 1294 13596 1300
rect 14568 1222 14596 3470
rect 14648 3120 14700 3126
rect 14648 3062 14700 3068
rect 14660 2854 14688 3062
rect 14936 2854 14964 5102
rect 15120 4486 15148 5170
rect 15212 5098 15240 7754
rect 15384 7336 15436 7342
rect 15384 7278 15436 7284
rect 15396 6914 15424 7278
rect 15580 6914 15608 11222
rect 15948 9081 15976 17546
rect 16040 16726 16068 17614
rect 16120 17536 16172 17542
rect 16120 17478 16172 17484
rect 16028 16720 16080 16726
rect 16028 16662 16080 16668
rect 16132 16572 16160 17478
rect 16214 17436 16522 17445
rect 16214 17434 16220 17436
rect 16276 17434 16300 17436
rect 16356 17434 16380 17436
rect 16436 17434 16460 17436
rect 16516 17434 16522 17436
rect 16276 17382 16278 17434
rect 16458 17382 16460 17434
rect 16214 17380 16220 17382
rect 16276 17380 16300 17382
rect 16356 17380 16380 17382
rect 16436 17380 16460 17382
rect 16516 17380 16522 17382
rect 16214 17371 16522 17380
rect 16948 17196 17000 17202
rect 16948 17138 17000 17144
rect 16580 16992 16632 16998
rect 16580 16934 16632 16940
rect 16212 16584 16264 16590
rect 16040 16544 16212 16572
rect 16040 13530 16068 16544
rect 16212 16526 16264 16532
rect 16214 16348 16522 16357
rect 16214 16346 16220 16348
rect 16276 16346 16300 16348
rect 16356 16346 16380 16348
rect 16436 16346 16460 16348
rect 16516 16346 16522 16348
rect 16276 16294 16278 16346
rect 16458 16294 16460 16346
rect 16214 16292 16220 16294
rect 16276 16292 16300 16294
rect 16356 16292 16380 16294
rect 16436 16292 16460 16294
rect 16516 16292 16522 16294
rect 16214 16283 16522 16292
rect 16212 16176 16264 16182
rect 16212 16118 16264 16124
rect 16224 15570 16252 16118
rect 16212 15564 16264 15570
rect 16212 15506 16264 15512
rect 16224 15450 16252 15506
rect 16592 15502 16620 16934
rect 16960 16726 16988 17138
rect 17132 17060 17184 17066
rect 17132 17002 17184 17008
rect 17040 16992 17092 16998
rect 17040 16934 17092 16940
rect 16948 16720 17000 16726
rect 16948 16662 17000 16668
rect 16764 16652 16816 16658
rect 16764 16594 16816 16600
rect 16776 16454 16804 16594
rect 16764 16448 16816 16454
rect 16764 16390 16816 16396
rect 16776 16114 16804 16390
rect 16960 16250 16988 16662
rect 16948 16244 17000 16250
rect 16948 16186 17000 16192
rect 17052 16153 17080 16934
rect 17144 16522 17172 17002
rect 17132 16516 17184 16522
rect 17132 16458 17184 16464
rect 17038 16144 17094 16153
rect 16764 16108 16816 16114
rect 17144 16114 17172 16458
rect 17038 16079 17094 16088
rect 17132 16108 17184 16114
rect 16764 16050 16816 16056
rect 17132 16050 17184 16056
rect 17328 15910 17356 21270
rect 17498 21200 17554 21270
rect 19522 21200 19578 22000
rect 21546 21200 21602 22000
rect 23570 21200 23626 22000
rect 25594 21200 25650 22000
rect 17592 19304 17644 19310
rect 17592 19246 17644 19252
rect 17604 18834 17632 19246
rect 17592 18828 17644 18834
rect 17592 18770 17644 18776
rect 17500 18760 17552 18766
rect 17500 18702 17552 18708
rect 17512 18086 17540 18702
rect 18144 18624 18196 18630
rect 18144 18566 18196 18572
rect 18156 18358 18184 18566
rect 18144 18352 18196 18358
rect 18144 18294 18196 18300
rect 17960 18148 18012 18154
rect 17960 18090 18012 18096
rect 17500 18080 17552 18086
rect 17500 18022 17552 18028
rect 17512 17542 17540 18022
rect 17972 17678 18000 18090
rect 17960 17672 18012 17678
rect 17960 17614 18012 17620
rect 18236 17604 18288 17610
rect 18236 17546 18288 17552
rect 17500 17536 17552 17542
rect 17500 17478 17552 17484
rect 18248 17202 18276 17546
rect 18420 17536 18472 17542
rect 18420 17478 18472 17484
rect 18236 17196 18288 17202
rect 18236 17138 18288 17144
rect 18248 16590 18276 17138
rect 18432 16726 18460 17478
rect 19340 17196 19392 17202
rect 19340 17138 19392 17144
rect 18420 16720 18472 16726
rect 18420 16662 18472 16668
rect 19352 16590 19380 17138
rect 19536 17066 19564 21200
rect 20214 20156 20522 20165
rect 20214 20154 20220 20156
rect 20276 20154 20300 20156
rect 20356 20154 20380 20156
rect 20436 20154 20460 20156
rect 20516 20154 20522 20156
rect 20276 20102 20278 20154
rect 20458 20102 20460 20154
rect 20214 20100 20220 20102
rect 20276 20100 20300 20102
rect 20356 20100 20380 20102
rect 20436 20100 20460 20102
rect 20516 20100 20522 20102
rect 20214 20091 20522 20100
rect 20214 19068 20522 19077
rect 20214 19066 20220 19068
rect 20276 19066 20300 19068
rect 20356 19066 20380 19068
rect 20436 19066 20460 19068
rect 20516 19066 20522 19068
rect 20276 19014 20278 19066
rect 20458 19014 20460 19066
rect 20214 19012 20220 19014
rect 20276 19012 20300 19014
rect 20356 19012 20380 19014
rect 20436 19012 20460 19014
rect 20516 19012 20522 19014
rect 20214 19003 20522 19012
rect 20214 17980 20522 17989
rect 20214 17978 20220 17980
rect 20276 17978 20300 17980
rect 20356 17978 20380 17980
rect 20436 17978 20460 17980
rect 20516 17978 20522 17980
rect 20276 17926 20278 17978
rect 20458 17926 20460 17978
rect 20214 17924 20220 17926
rect 20276 17924 20300 17926
rect 20356 17924 20380 17926
rect 20436 17924 20460 17926
rect 20516 17924 20522 17926
rect 20214 17915 20522 17924
rect 19524 17060 19576 17066
rect 19524 17002 19576 17008
rect 21560 16998 21588 21200
rect 21548 16992 21600 16998
rect 21548 16934 21600 16940
rect 20214 16892 20522 16901
rect 20214 16890 20220 16892
rect 20276 16890 20300 16892
rect 20356 16890 20380 16892
rect 20436 16890 20460 16892
rect 20516 16890 20522 16892
rect 20276 16838 20278 16890
rect 20458 16838 20460 16890
rect 20214 16836 20220 16838
rect 20276 16836 20300 16838
rect 20356 16836 20380 16838
rect 20436 16836 20460 16838
rect 20516 16836 20522 16838
rect 20214 16827 20522 16836
rect 23584 16794 23612 21200
rect 24214 20700 24522 20709
rect 24214 20698 24220 20700
rect 24276 20698 24300 20700
rect 24356 20698 24380 20700
rect 24436 20698 24460 20700
rect 24516 20698 24522 20700
rect 24276 20646 24278 20698
rect 24458 20646 24460 20698
rect 24214 20644 24220 20646
rect 24276 20644 24300 20646
rect 24356 20644 24380 20646
rect 24436 20644 24460 20646
rect 24516 20644 24522 20646
rect 24214 20635 24522 20644
rect 24860 19984 24912 19990
rect 24860 19926 24912 19932
rect 24872 19689 24900 19926
rect 24858 19680 24914 19689
rect 24214 19612 24522 19621
rect 24858 19615 24914 19624
rect 24214 19610 24220 19612
rect 24276 19610 24300 19612
rect 24356 19610 24380 19612
rect 24436 19610 24460 19612
rect 24516 19610 24522 19612
rect 24276 19558 24278 19610
rect 24458 19558 24460 19610
rect 24214 19556 24220 19558
rect 24276 19556 24300 19558
rect 24356 19556 24380 19558
rect 24436 19556 24460 19558
rect 24516 19556 24522 19558
rect 24214 19547 24522 19556
rect 25608 19310 25636 21200
rect 25596 19304 25648 19310
rect 25596 19246 25648 19252
rect 24952 19168 25004 19174
rect 24952 19110 25004 19116
rect 24214 18524 24522 18533
rect 24214 18522 24220 18524
rect 24276 18522 24300 18524
rect 24356 18522 24380 18524
rect 24436 18522 24460 18524
rect 24516 18522 24522 18524
rect 24276 18470 24278 18522
rect 24458 18470 24460 18522
rect 24214 18468 24220 18470
rect 24276 18468 24300 18470
rect 24356 18468 24380 18470
rect 24436 18468 24460 18470
rect 24516 18468 24522 18470
rect 24214 18459 24522 18468
rect 24860 18420 24912 18426
rect 24860 18362 24912 18368
rect 24214 17436 24522 17445
rect 24214 17434 24220 17436
rect 24276 17434 24300 17436
rect 24356 17434 24380 17436
rect 24436 17434 24460 17436
rect 24516 17434 24522 17436
rect 24276 17382 24278 17434
rect 24458 17382 24460 17434
rect 24214 17380 24220 17382
rect 24276 17380 24300 17382
rect 24356 17380 24380 17382
rect 24436 17380 24460 17382
rect 24516 17380 24522 17382
rect 24214 17371 24522 17380
rect 23572 16788 23624 16794
rect 23572 16730 23624 16736
rect 18236 16584 18288 16590
rect 18236 16526 18288 16532
rect 19340 16584 19392 16590
rect 19340 16526 19392 16532
rect 24214 16348 24522 16357
rect 24214 16346 24220 16348
rect 24276 16346 24300 16348
rect 24356 16346 24380 16348
rect 24436 16346 24460 16348
rect 24516 16346 24522 16348
rect 24276 16294 24278 16346
rect 24458 16294 24460 16346
rect 24214 16292 24220 16294
rect 24276 16292 24300 16294
rect 24356 16292 24380 16294
rect 24436 16292 24460 16294
rect 24516 16292 24522 16294
rect 24214 16283 24522 16292
rect 24872 16153 24900 18362
rect 24858 16144 24914 16153
rect 24858 16079 24914 16088
rect 17316 15904 17368 15910
rect 17316 15846 17368 15852
rect 20214 15804 20522 15813
rect 20214 15802 20220 15804
rect 20276 15802 20300 15804
rect 20356 15802 20380 15804
rect 20436 15802 20460 15804
rect 20516 15802 20522 15804
rect 20276 15750 20278 15802
rect 20458 15750 20460 15802
rect 20214 15748 20220 15750
rect 20276 15748 20300 15750
rect 20356 15748 20380 15750
rect 20436 15748 20460 15750
rect 20516 15748 20522 15750
rect 20214 15739 20522 15748
rect 16132 15422 16252 15450
rect 16580 15496 16632 15502
rect 16580 15438 16632 15444
rect 16132 15094 16160 15422
rect 16214 15260 16522 15269
rect 16214 15258 16220 15260
rect 16276 15258 16300 15260
rect 16356 15258 16380 15260
rect 16436 15258 16460 15260
rect 16516 15258 16522 15260
rect 16276 15206 16278 15258
rect 16458 15206 16460 15258
rect 16214 15204 16220 15206
rect 16276 15204 16300 15206
rect 16356 15204 16380 15206
rect 16436 15204 16460 15206
rect 16516 15204 16522 15206
rect 16214 15195 16522 15204
rect 24214 15260 24522 15269
rect 24214 15258 24220 15260
rect 24276 15258 24300 15260
rect 24356 15258 24380 15260
rect 24436 15258 24460 15260
rect 24516 15258 24522 15260
rect 24276 15206 24278 15258
rect 24458 15206 24460 15258
rect 24214 15204 24220 15206
rect 24276 15204 24300 15206
rect 24356 15204 24380 15206
rect 24436 15204 24460 15206
rect 24516 15204 24522 15206
rect 24214 15195 24522 15204
rect 16120 15088 16172 15094
rect 16120 15030 16172 15036
rect 16132 14414 16160 15030
rect 16304 15020 16356 15026
rect 16304 14962 16356 14968
rect 16948 15020 17000 15026
rect 16948 14962 17000 14968
rect 16316 14482 16344 14962
rect 16856 14816 16908 14822
rect 16856 14758 16908 14764
rect 16304 14476 16356 14482
rect 16304 14418 16356 14424
rect 16120 14408 16172 14414
rect 16120 14350 16172 14356
rect 16214 14172 16522 14181
rect 16214 14170 16220 14172
rect 16276 14170 16300 14172
rect 16356 14170 16380 14172
rect 16436 14170 16460 14172
rect 16516 14170 16522 14172
rect 16276 14118 16278 14170
rect 16458 14118 16460 14170
rect 16214 14116 16220 14118
rect 16276 14116 16300 14118
rect 16356 14116 16380 14118
rect 16436 14116 16460 14118
rect 16516 14116 16522 14118
rect 16214 14107 16522 14116
rect 16868 14074 16896 14758
rect 16960 14618 16988 14962
rect 20214 14716 20522 14725
rect 20214 14714 20220 14716
rect 20276 14714 20300 14716
rect 20356 14714 20380 14716
rect 20436 14714 20460 14716
rect 20516 14714 20522 14716
rect 20276 14662 20278 14714
rect 20458 14662 20460 14714
rect 20214 14660 20220 14662
rect 20276 14660 20300 14662
rect 20356 14660 20380 14662
rect 20436 14660 20460 14662
rect 20516 14660 20522 14662
rect 20214 14651 20522 14660
rect 16948 14612 17000 14618
rect 16948 14554 17000 14560
rect 24214 14172 24522 14181
rect 24214 14170 24220 14172
rect 24276 14170 24300 14172
rect 24356 14170 24380 14172
rect 24436 14170 24460 14172
rect 24516 14170 24522 14172
rect 24276 14118 24278 14170
rect 24458 14118 24460 14170
rect 24214 14116 24220 14118
rect 24276 14116 24300 14118
rect 24356 14116 24380 14118
rect 24436 14116 24460 14118
rect 24516 14116 24522 14118
rect 24214 14107 24522 14116
rect 16856 14068 16908 14074
rect 16856 14010 16908 14016
rect 16764 13932 16816 13938
rect 16764 13874 16816 13880
rect 16028 13524 16080 13530
rect 16028 13466 16080 13472
rect 16040 12918 16068 13466
rect 16776 13326 16804 13874
rect 16764 13320 16816 13326
rect 16764 13262 16816 13268
rect 16214 13084 16522 13093
rect 16214 13082 16220 13084
rect 16276 13082 16300 13084
rect 16356 13082 16380 13084
rect 16436 13082 16460 13084
rect 16516 13082 16522 13084
rect 16276 13030 16278 13082
rect 16458 13030 16460 13082
rect 16214 13028 16220 13030
rect 16276 13028 16300 13030
rect 16356 13028 16380 13030
rect 16436 13028 16460 13030
rect 16516 13028 16522 13030
rect 16214 13019 16522 13028
rect 16028 12912 16080 12918
rect 16028 12854 16080 12860
rect 16672 12640 16724 12646
rect 16672 12582 16724 12588
rect 16580 12096 16632 12102
rect 16580 12038 16632 12044
rect 16214 11996 16522 12005
rect 16214 11994 16220 11996
rect 16276 11994 16300 11996
rect 16356 11994 16380 11996
rect 16436 11994 16460 11996
rect 16516 11994 16522 11996
rect 16276 11942 16278 11994
rect 16458 11942 16460 11994
rect 16214 11940 16220 11942
rect 16276 11940 16300 11942
rect 16356 11940 16380 11942
rect 16436 11940 16460 11942
rect 16516 11940 16522 11942
rect 16214 11931 16522 11940
rect 16592 11762 16620 12038
rect 16580 11756 16632 11762
rect 16580 11698 16632 11704
rect 16028 11620 16080 11626
rect 16028 11562 16080 11568
rect 16040 10538 16068 11562
rect 16214 10908 16522 10917
rect 16214 10906 16220 10908
rect 16276 10906 16300 10908
rect 16356 10906 16380 10908
rect 16436 10906 16460 10908
rect 16516 10906 16522 10908
rect 16276 10854 16278 10906
rect 16458 10854 16460 10906
rect 16214 10852 16220 10854
rect 16276 10852 16300 10854
rect 16356 10852 16380 10854
rect 16436 10852 16460 10854
rect 16516 10852 16522 10854
rect 16214 10843 16522 10852
rect 16120 10668 16172 10674
rect 16120 10610 16172 10616
rect 16028 10532 16080 10538
rect 16028 10474 16080 10480
rect 16040 10062 16068 10474
rect 16132 10062 16160 10610
rect 16592 10130 16620 11698
rect 16684 11082 16712 12582
rect 16776 12442 16804 13262
rect 16764 12436 16816 12442
rect 16764 12378 16816 12384
rect 16868 12306 16896 14010
rect 20214 13628 20522 13637
rect 20214 13626 20220 13628
rect 20276 13626 20300 13628
rect 20356 13626 20380 13628
rect 20436 13626 20460 13628
rect 20516 13626 20522 13628
rect 20276 13574 20278 13626
rect 20458 13574 20460 13626
rect 20214 13572 20220 13574
rect 20276 13572 20300 13574
rect 20356 13572 20380 13574
rect 20436 13572 20460 13574
rect 20516 13572 20522 13574
rect 20214 13563 20522 13572
rect 24214 13084 24522 13093
rect 24214 13082 24220 13084
rect 24276 13082 24300 13084
rect 24356 13082 24380 13084
rect 24436 13082 24460 13084
rect 24516 13082 24522 13084
rect 24276 13030 24278 13082
rect 24458 13030 24460 13082
rect 24214 13028 24220 13030
rect 24276 13028 24300 13030
rect 24356 13028 24380 13030
rect 24436 13028 24460 13030
rect 24516 13028 24522 13030
rect 24214 13019 24522 13028
rect 17868 12844 17920 12850
rect 17868 12786 17920 12792
rect 16948 12640 17000 12646
rect 16948 12582 17000 12588
rect 16764 12300 16816 12306
rect 16764 12242 16816 12248
rect 16856 12300 16908 12306
rect 16856 12242 16908 12248
rect 16776 12186 16804 12242
rect 16776 12158 16896 12186
rect 16960 12170 16988 12582
rect 17500 12300 17552 12306
rect 17500 12242 17552 12248
rect 16868 12102 16896 12158
rect 16948 12164 17000 12170
rect 16948 12106 17000 12112
rect 17224 12164 17276 12170
rect 17224 12106 17276 12112
rect 16856 12096 16908 12102
rect 16856 12038 16908 12044
rect 17236 11898 17264 12106
rect 17224 11892 17276 11898
rect 17224 11834 17276 11840
rect 17512 11762 17540 12242
rect 17880 12170 17908 12786
rect 24964 12617 24992 19110
rect 26148 16516 26200 16522
rect 26148 16458 26200 16464
rect 24950 12608 25006 12617
rect 20214 12540 20522 12549
rect 24950 12543 25006 12552
rect 20214 12538 20220 12540
rect 20276 12538 20300 12540
rect 20356 12538 20380 12540
rect 20436 12538 20460 12540
rect 20516 12538 20522 12540
rect 20276 12486 20278 12538
rect 20458 12486 20460 12538
rect 20214 12484 20220 12486
rect 20276 12484 20300 12486
rect 20356 12484 20380 12486
rect 20436 12484 20460 12486
rect 20516 12484 20522 12486
rect 20214 12475 20522 12484
rect 18236 12436 18288 12442
rect 18236 12378 18288 12384
rect 18248 12238 18276 12378
rect 19616 12300 19668 12306
rect 19616 12242 19668 12248
rect 18236 12232 18288 12238
rect 18512 12232 18564 12238
rect 18288 12180 18512 12186
rect 18236 12174 18564 12180
rect 17868 12164 17920 12170
rect 18248 12158 18552 12174
rect 19524 12164 19576 12170
rect 17868 12106 17920 12112
rect 19524 12106 19576 12112
rect 18328 12096 18380 12102
rect 18328 12038 18380 12044
rect 18340 11830 18368 12038
rect 18328 11824 18380 11830
rect 18328 11766 18380 11772
rect 16764 11756 16816 11762
rect 16764 11698 16816 11704
rect 17500 11756 17552 11762
rect 17500 11698 17552 11704
rect 16672 11076 16724 11082
rect 16672 11018 16724 11024
rect 16776 10810 16804 11698
rect 16948 11552 17000 11558
rect 16948 11494 17000 11500
rect 16960 11218 16988 11494
rect 17512 11218 17540 11698
rect 18052 11688 18104 11694
rect 18052 11630 18104 11636
rect 18064 11354 18092 11630
rect 19064 11620 19116 11626
rect 19064 11562 19116 11568
rect 18052 11348 18104 11354
rect 18052 11290 18104 11296
rect 16948 11212 17000 11218
rect 16948 11154 17000 11160
rect 17500 11212 17552 11218
rect 17500 11154 17552 11160
rect 16764 10804 16816 10810
rect 16764 10746 16816 10752
rect 17512 10674 17540 11154
rect 19076 11150 19104 11562
rect 19536 11354 19564 12106
rect 19524 11348 19576 11354
rect 19524 11290 19576 11296
rect 19064 11144 19116 11150
rect 19064 11086 19116 11092
rect 18052 11076 18104 11082
rect 18052 11018 18104 11024
rect 18064 10742 18092 11018
rect 18236 11008 18288 11014
rect 18236 10950 18288 10956
rect 18052 10736 18104 10742
rect 18052 10678 18104 10684
rect 16764 10668 16816 10674
rect 16764 10610 16816 10616
rect 17500 10668 17552 10674
rect 17500 10610 17552 10616
rect 16776 10266 16804 10610
rect 16948 10464 17000 10470
rect 16948 10406 17000 10412
rect 16764 10260 16816 10266
rect 16764 10202 16816 10208
rect 16580 10124 16632 10130
rect 16580 10066 16632 10072
rect 16028 10056 16080 10062
rect 16028 9998 16080 10004
rect 16120 10056 16172 10062
rect 16120 9998 16172 10004
rect 16214 9820 16522 9829
rect 16214 9818 16220 9820
rect 16276 9818 16300 9820
rect 16356 9818 16380 9820
rect 16436 9818 16460 9820
rect 16516 9818 16522 9820
rect 16276 9766 16278 9818
rect 16458 9766 16460 9818
rect 16214 9764 16220 9766
rect 16276 9764 16300 9766
rect 16356 9764 16380 9766
rect 16436 9764 16460 9766
rect 16516 9764 16522 9766
rect 16214 9755 16522 9764
rect 16960 9654 16988 10406
rect 18248 10130 18276 10950
rect 19156 10668 19208 10674
rect 19156 10610 19208 10616
rect 18788 10600 18840 10606
rect 18788 10542 18840 10548
rect 18696 10464 18748 10470
rect 18696 10406 18748 10412
rect 18236 10124 18288 10130
rect 18236 10066 18288 10072
rect 18708 10062 18736 10406
rect 18696 10056 18748 10062
rect 18696 9998 18748 10004
rect 17776 9988 17828 9994
rect 17776 9930 17828 9936
rect 16948 9648 17000 9654
rect 16948 9590 17000 9596
rect 17684 9648 17736 9654
rect 17684 9590 17736 9596
rect 16672 9512 16724 9518
rect 16672 9454 16724 9460
rect 15934 9072 15990 9081
rect 15934 9007 15990 9016
rect 15660 8968 15712 8974
rect 15660 8910 15712 8916
rect 16488 8968 16540 8974
rect 16488 8910 16540 8916
rect 15672 7886 15700 8910
rect 16028 8900 16080 8906
rect 16028 8842 16080 8848
rect 16040 7886 16068 8842
rect 16500 8838 16528 8910
rect 16488 8832 16540 8838
rect 16488 8774 16540 8780
rect 16214 8732 16522 8741
rect 16214 8730 16220 8732
rect 16276 8730 16300 8732
rect 16356 8730 16380 8732
rect 16436 8730 16460 8732
rect 16516 8730 16522 8732
rect 16276 8678 16278 8730
rect 16458 8678 16460 8730
rect 16214 8676 16220 8678
rect 16276 8676 16300 8678
rect 16356 8676 16380 8678
rect 16436 8676 16460 8678
rect 16516 8676 16522 8678
rect 16214 8667 16522 8676
rect 16684 8430 16712 9454
rect 17696 9178 17724 9590
rect 17788 9518 17816 9930
rect 17776 9512 17828 9518
rect 17776 9454 17828 9460
rect 17684 9172 17736 9178
rect 17684 9114 17736 9120
rect 17224 9104 17276 9110
rect 17224 9046 17276 9052
rect 17236 8634 17264 9046
rect 17500 8900 17552 8906
rect 17500 8842 17552 8848
rect 17224 8628 17276 8634
rect 17224 8570 17276 8576
rect 17512 8430 17540 8842
rect 17788 8634 17816 9454
rect 18420 9376 18472 9382
rect 18420 9318 18472 9324
rect 18432 9042 18460 9318
rect 18420 9036 18472 9042
rect 18420 8978 18472 8984
rect 17960 8968 18012 8974
rect 17960 8910 18012 8916
rect 17776 8628 17828 8634
rect 17776 8570 17828 8576
rect 17592 8492 17644 8498
rect 17592 8434 17644 8440
rect 16672 8424 16724 8430
rect 16672 8366 16724 8372
rect 17500 8424 17552 8430
rect 17500 8366 17552 8372
rect 16684 7886 16712 8366
rect 16948 8288 17000 8294
rect 16948 8230 17000 8236
rect 16960 7954 16988 8230
rect 16948 7948 17000 7954
rect 16948 7890 17000 7896
rect 15660 7880 15712 7886
rect 15660 7822 15712 7828
rect 16028 7880 16080 7886
rect 16028 7822 16080 7828
rect 16672 7880 16724 7886
rect 16672 7822 16724 7828
rect 15672 7410 15700 7822
rect 15844 7744 15896 7750
rect 15844 7686 15896 7692
rect 15660 7404 15712 7410
rect 15660 7346 15712 7352
rect 15396 6886 15516 6914
rect 15580 6886 15700 6914
rect 15488 6662 15516 6886
rect 15672 6798 15700 6886
rect 15660 6792 15712 6798
rect 15660 6734 15712 6740
rect 15476 6656 15528 6662
rect 15476 6598 15528 6604
rect 15488 5302 15516 6598
rect 15856 6322 15884 7686
rect 16214 7644 16522 7653
rect 16214 7642 16220 7644
rect 16276 7642 16300 7644
rect 16356 7642 16380 7644
rect 16436 7642 16460 7644
rect 16516 7642 16522 7644
rect 16276 7590 16278 7642
rect 16458 7590 16460 7642
rect 16214 7588 16220 7590
rect 16276 7588 16300 7590
rect 16356 7588 16380 7590
rect 16436 7588 16460 7590
rect 16516 7588 16522 7590
rect 16214 7579 16522 7588
rect 16684 7546 16712 7822
rect 17604 7750 17632 8434
rect 17592 7744 17644 7750
rect 17592 7686 17644 7692
rect 16672 7540 16724 7546
rect 16672 7482 16724 7488
rect 16214 6556 16522 6565
rect 16214 6554 16220 6556
rect 16276 6554 16300 6556
rect 16356 6554 16380 6556
rect 16436 6554 16460 6556
rect 16516 6554 16522 6556
rect 16276 6502 16278 6554
rect 16458 6502 16460 6554
rect 16214 6500 16220 6502
rect 16276 6500 16300 6502
rect 16356 6500 16380 6502
rect 16436 6500 16460 6502
rect 16516 6500 16522 6502
rect 16214 6491 16522 6500
rect 15844 6316 15896 6322
rect 15844 6258 15896 6264
rect 15936 6112 15988 6118
rect 15936 6054 15988 6060
rect 15750 5672 15806 5681
rect 15750 5607 15806 5616
rect 15764 5370 15792 5607
rect 15948 5574 15976 6054
rect 16120 5772 16172 5778
rect 16120 5714 16172 5720
rect 15936 5568 15988 5574
rect 15936 5510 15988 5516
rect 16132 5370 16160 5714
rect 16684 5642 16712 7482
rect 16948 7404 17000 7410
rect 16948 7346 17000 7352
rect 16960 6322 16988 7346
rect 17132 6860 17184 6866
rect 17132 6802 17184 6808
rect 16948 6316 17000 6322
rect 16948 6258 17000 6264
rect 16672 5636 16724 5642
rect 16672 5578 16724 5584
rect 16214 5468 16522 5477
rect 16214 5466 16220 5468
rect 16276 5466 16300 5468
rect 16356 5466 16380 5468
rect 16436 5466 16460 5468
rect 16516 5466 16522 5468
rect 16276 5414 16278 5466
rect 16458 5414 16460 5466
rect 16214 5412 16220 5414
rect 16276 5412 16300 5414
rect 16356 5412 16380 5414
rect 16436 5412 16460 5414
rect 16516 5412 16522 5414
rect 16214 5403 16522 5412
rect 15752 5364 15804 5370
rect 15752 5306 15804 5312
rect 16120 5364 16172 5370
rect 16120 5306 16172 5312
rect 15476 5296 15528 5302
rect 15476 5238 15528 5244
rect 16028 5228 16080 5234
rect 16028 5170 16080 5176
rect 16120 5228 16172 5234
rect 16120 5170 16172 5176
rect 15200 5092 15252 5098
rect 15200 5034 15252 5040
rect 15844 5092 15896 5098
rect 15844 5034 15896 5040
rect 15108 4480 15160 4486
rect 15108 4422 15160 4428
rect 15016 3392 15068 3398
rect 15016 3334 15068 3340
rect 14648 2848 14700 2854
rect 14648 2790 14700 2796
rect 14924 2848 14976 2854
rect 14924 2790 14976 2796
rect 14936 1494 14964 2790
rect 15028 2038 15056 3334
rect 15016 2032 15068 2038
rect 15016 1974 15068 1980
rect 14924 1488 14976 1494
rect 14924 1430 14976 1436
rect 15120 1290 15148 4422
rect 15856 3058 15884 5034
rect 16040 4758 16068 5170
rect 16028 4752 16080 4758
rect 16028 4694 16080 4700
rect 16040 4010 16068 4694
rect 16132 4554 16160 5170
rect 16120 4548 16172 4554
rect 16120 4490 16172 4496
rect 16132 4078 16160 4490
rect 16214 4380 16522 4389
rect 16214 4378 16220 4380
rect 16276 4378 16300 4380
rect 16356 4378 16380 4380
rect 16436 4378 16460 4380
rect 16516 4378 16522 4380
rect 16276 4326 16278 4378
rect 16458 4326 16460 4378
rect 16214 4324 16220 4326
rect 16276 4324 16300 4326
rect 16356 4324 16380 4326
rect 16436 4324 16460 4326
rect 16516 4324 16522 4326
rect 16214 4315 16522 4324
rect 16488 4208 16540 4214
rect 16488 4150 16540 4156
rect 16120 4072 16172 4078
rect 16120 4014 16172 4020
rect 16028 4004 16080 4010
rect 16028 3946 16080 3952
rect 16500 3738 16528 4150
rect 16684 4010 16712 5578
rect 16960 5234 16988 6258
rect 17040 6112 17092 6118
rect 17040 6054 17092 6060
rect 16948 5228 17000 5234
rect 16948 5170 17000 5176
rect 16960 4826 16988 5170
rect 17052 5166 17080 6054
rect 17040 5160 17092 5166
rect 17040 5102 17092 5108
rect 16948 4820 17000 4826
rect 16948 4762 17000 4768
rect 16672 4004 16724 4010
rect 16672 3946 16724 3952
rect 16488 3732 16540 3738
rect 16488 3674 16540 3680
rect 16684 3670 16712 3946
rect 16672 3664 16724 3670
rect 16672 3606 16724 3612
rect 15936 3596 15988 3602
rect 15936 3538 15988 3544
rect 15660 3052 15712 3058
rect 15660 2994 15712 3000
rect 15844 3052 15896 3058
rect 15844 2994 15896 3000
rect 15672 2514 15700 2994
rect 15948 2514 15976 3538
rect 16672 3528 16724 3534
rect 16672 3470 16724 3476
rect 16214 3292 16522 3301
rect 16214 3290 16220 3292
rect 16276 3290 16300 3292
rect 16356 3290 16380 3292
rect 16436 3290 16460 3292
rect 16516 3290 16522 3292
rect 16276 3238 16278 3290
rect 16458 3238 16460 3290
rect 16214 3236 16220 3238
rect 16276 3236 16300 3238
rect 16356 3236 16380 3238
rect 16436 3236 16460 3238
rect 16516 3236 16522 3238
rect 16214 3227 16522 3236
rect 16212 3188 16264 3194
rect 16212 3130 16264 3136
rect 16224 2650 16252 3130
rect 16684 3058 16712 3470
rect 16672 3052 16724 3058
rect 16672 2994 16724 3000
rect 16948 2984 17000 2990
rect 16948 2926 17000 2932
rect 16580 2848 16632 2854
rect 16580 2790 16632 2796
rect 16960 2802 16988 2926
rect 17052 2922 17080 5102
rect 17144 4826 17172 6802
rect 17224 6112 17276 6118
rect 17224 6054 17276 6060
rect 17236 5642 17264 6054
rect 17224 5636 17276 5642
rect 17224 5578 17276 5584
rect 17132 4820 17184 4826
rect 17132 4762 17184 4768
rect 17144 4078 17172 4762
rect 17500 4480 17552 4486
rect 17500 4422 17552 4428
rect 17132 4072 17184 4078
rect 17132 4014 17184 4020
rect 17512 3602 17540 4422
rect 17604 4282 17632 7686
rect 17776 7404 17828 7410
rect 17776 7346 17828 7352
rect 17788 6662 17816 7346
rect 17972 6934 18000 8910
rect 18708 8634 18736 9998
rect 18800 9722 18828 10542
rect 19168 10266 19196 10610
rect 19628 10606 19656 12242
rect 20996 12096 21048 12102
rect 20996 12038 21048 12044
rect 21008 11762 21036 12038
rect 24214 11996 24522 12005
rect 24214 11994 24220 11996
rect 24276 11994 24300 11996
rect 24356 11994 24380 11996
rect 24436 11994 24460 11996
rect 24516 11994 24522 11996
rect 24276 11942 24278 11994
rect 24458 11942 24460 11994
rect 24214 11940 24220 11942
rect 24276 11940 24300 11942
rect 24356 11940 24380 11942
rect 24436 11940 24460 11942
rect 24516 11940 24522 11942
rect 24214 11931 24522 11940
rect 20996 11756 21048 11762
rect 20996 11698 21048 11704
rect 19984 11688 20036 11694
rect 19984 11630 20036 11636
rect 19800 11552 19852 11558
rect 19800 11494 19852 11500
rect 19812 11150 19840 11494
rect 19996 11218 20024 11630
rect 20214 11452 20522 11461
rect 20214 11450 20220 11452
rect 20276 11450 20300 11452
rect 20356 11450 20380 11452
rect 20436 11450 20460 11452
rect 20516 11450 20522 11452
rect 20276 11398 20278 11450
rect 20458 11398 20460 11450
rect 20214 11396 20220 11398
rect 20276 11396 20300 11398
rect 20356 11396 20380 11398
rect 20436 11396 20460 11398
rect 20516 11396 20522 11398
rect 20214 11387 20522 11396
rect 21008 11218 21036 11698
rect 22652 11620 22704 11626
rect 22652 11562 22704 11568
rect 22284 11348 22336 11354
rect 22284 11290 22336 11296
rect 19984 11212 20036 11218
rect 19984 11154 20036 11160
rect 20996 11212 21048 11218
rect 20996 11154 21048 11160
rect 19800 11144 19852 11150
rect 19800 11086 19852 11092
rect 19616 10600 19668 10606
rect 19616 10542 19668 10548
rect 19156 10260 19208 10266
rect 19156 10202 19208 10208
rect 19628 10130 19656 10542
rect 19616 10124 19668 10130
rect 19616 10066 19668 10072
rect 19156 10056 19208 10062
rect 19524 10056 19576 10062
rect 19156 9998 19208 10004
rect 19260 10016 19524 10044
rect 18972 9920 19024 9926
rect 18972 9862 19024 9868
rect 18788 9716 18840 9722
rect 18788 9658 18840 9664
rect 18984 9586 19012 9862
rect 18972 9580 19024 9586
rect 18972 9522 19024 9528
rect 19168 8906 19196 9998
rect 19156 8900 19208 8906
rect 19156 8842 19208 8848
rect 18696 8628 18748 8634
rect 18696 8570 18748 8576
rect 19260 8566 19288 10016
rect 19524 9998 19576 10004
rect 19628 9874 19656 10066
rect 19536 9846 19656 9874
rect 19536 9722 19564 9846
rect 19524 9716 19576 9722
rect 19524 9658 19576 9664
rect 19536 9586 19564 9658
rect 19524 9580 19576 9586
rect 19524 9522 19576 9528
rect 19800 9512 19852 9518
rect 19800 9454 19852 9460
rect 19524 8832 19576 8838
rect 19524 8774 19576 8780
rect 18972 8560 19024 8566
rect 18972 8502 19024 8508
rect 19248 8560 19300 8566
rect 19248 8502 19300 8508
rect 18788 8492 18840 8498
rect 18788 8434 18840 8440
rect 18236 8084 18288 8090
rect 18236 8026 18288 8032
rect 17960 6928 18012 6934
rect 17960 6870 18012 6876
rect 17972 6798 18000 6870
rect 18248 6798 18276 8026
rect 18800 7342 18828 8434
rect 18984 7886 19012 8502
rect 19536 8498 19564 8774
rect 19812 8634 19840 9454
rect 19996 9042 20024 11154
rect 20076 11008 20128 11014
rect 20076 10950 20128 10956
rect 21916 11008 21968 11014
rect 21916 10950 21968 10956
rect 20088 9994 20116 10950
rect 21180 10668 21232 10674
rect 21100 10628 21180 10656
rect 20214 10364 20522 10373
rect 20214 10362 20220 10364
rect 20276 10362 20300 10364
rect 20356 10362 20380 10364
rect 20436 10362 20460 10364
rect 20516 10362 20522 10364
rect 20276 10310 20278 10362
rect 20458 10310 20460 10362
rect 20214 10308 20220 10310
rect 20276 10308 20300 10310
rect 20356 10308 20380 10310
rect 20436 10308 20460 10310
rect 20516 10308 20522 10310
rect 20214 10299 20522 10308
rect 21100 10130 21128 10628
rect 21180 10610 21232 10616
rect 21732 10668 21784 10674
rect 21732 10610 21784 10616
rect 21180 10464 21232 10470
rect 21180 10406 21232 10412
rect 21088 10124 21140 10130
rect 21088 10066 21140 10072
rect 21192 9994 21220 10406
rect 21456 10124 21508 10130
rect 21456 10066 21508 10072
rect 20076 9988 20128 9994
rect 20076 9930 20128 9936
rect 21180 9988 21232 9994
rect 21180 9930 21232 9936
rect 20904 9580 20956 9586
rect 20904 9522 20956 9528
rect 20214 9276 20522 9285
rect 20214 9274 20220 9276
rect 20276 9274 20300 9276
rect 20356 9274 20380 9276
rect 20436 9274 20460 9276
rect 20516 9274 20522 9276
rect 20276 9222 20278 9274
rect 20458 9222 20460 9274
rect 20214 9220 20220 9222
rect 20276 9220 20300 9222
rect 20356 9220 20380 9222
rect 20436 9220 20460 9222
rect 20516 9220 20522 9222
rect 20214 9211 20522 9220
rect 19984 9036 20036 9042
rect 19984 8978 20036 8984
rect 19800 8628 19852 8634
rect 19800 8570 19852 8576
rect 19524 8492 19576 8498
rect 19524 8434 19576 8440
rect 19616 8424 19668 8430
rect 19616 8366 19668 8372
rect 19432 8356 19484 8362
rect 19432 8298 19484 8304
rect 19444 7886 19472 8298
rect 18972 7880 19024 7886
rect 18972 7822 19024 7828
rect 19432 7880 19484 7886
rect 19432 7822 19484 7828
rect 18880 7744 18932 7750
rect 18880 7686 18932 7692
rect 18892 7478 18920 7686
rect 18880 7472 18932 7478
rect 18880 7414 18932 7420
rect 18788 7336 18840 7342
rect 18788 7278 18840 7284
rect 18604 6996 18656 7002
rect 18604 6938 18656 6944
rect 17960 6792 18012 6798
rect 17960 6734 18012 6740
rect 18236 6792 18288 6798
rect 18236 6734 18288 6740
rect 17776 6656 17828 6662
rect 17776 6598 17828 6604
rect 18616 6322 18644 6938
rect 17684 6316 17736 6322
rect 17684 6258 17736 6264
rect 18604 6316 18656 6322
rect 18604 6258 18656 6264
rect 17696 5370 17724 6258
rect 18236 6112 18288 6118
rect 18236 6054 18288 6060
rect 18248 5642 18276 6054
rect 18236 5636 18288 5642
rect 18236 5578 18288 5584
rect 18144 5568 18196 5574
rect 18144 5510 18196 5516
rect 18156 5370 18184 5510
rect 17684 5364 17736 5370
rect 17684 5306 17736 5312
rect 18144 5364 18196 5370
rect 18144 5306 18196 5312
rect 18800 4690 18828 7278
rect 18984 6934 19012 7822
rect 19432 7472 19484 7478
rect 19432 7414 19484 7420
rect 19248 7404 19300 7410
rect 19248 7346 19300 7352
rect 19260 7002 19288 7346
rect 19248 6996 19300 7002
rect 19248 6938 19300 6944
rect 18972 6928 19024 6934
rect 18972 6870 19024 6876
rect 19156 6316 19208 6322
rect 19156 6258 19208 6264
rect 19168 5234 19196 6258
rect 19444 5914 19472 7414
rect 19524 6996 19576 7002
rect 19524 6938 19576 6944
rect 19536 6798 19564 6938
rect 19524 6792 19576 6798
rect 19524 6734 19576 6740
rect 19432 5908 19484 5914
rect 19432 5850 19484 5856
rect 19536 5778 19564 6734
rect 19628 6254 19656 8366
rect 19616 6248 19668 6254
rect 19616 6190 19668 6196
rect 19524 5772 19576 5778
rect 19524 5714 19576 5720
rect 19156 5228 19208 5234
rect 19156 5170 19208 5176
rect 19340 4752 19392 4758
rect 19340 4694 19392 4700
rect 18788 4684 18840 4690
rect 18788 4626 18840 4632
rect 17684 4616 17736 4622
rect 17684 4558 17736 4564
rect 17696 4282 17724 4558
rect 18512 4480 18564 4486
rect 18512 4422 18564 4428
rect 17592 4276 17644 4282
rect 17592 4218 17644 4224
rect 17684 4276 17736 4282
rect 17684 4218 17736 4224
rect 18524 4214 18552 4422
rect 19352 4282 19380 4694
rect 19340 4276 19392 4282
rect 19340 4218 19392 4224
rect 18512 4208 18564 4214
rect 18512 4150 18564 4156
rect 17592 4072 17644 4078
rect 17592 4014 17644 4020
rect 17604 3738 17632 4014
rect 18052 3936 18104 3942
rect 18052 3878 18104 3884
rect 17592 3732 17644 3738
rect 17592 3674 17644 3680
rect 17500 3596 17552 3602
rect 17500 3538 17552 3544
rect 17604 3194 17632 3674
rect 18064 3602 18092 3878
rect 18052 3596 18104 3602
rect 18052 3538 18104 3544
rect 19352 3534 19380 4218
rect 19628 4010 19656 6190
rect 19708 6112 19760 6118
rect 19708 6054 19760 6060
rect 19800 6112 19852 6118
rect 19800 6054 19852 6060
rect 19720 5302 19748 6054
rect 19812 5778 19840 6054
rect 19800 5772 19852 5778
rect 19800 5714 19852 5720
rect 19708 5296 19760 5302
rect 19708 5238 19760 5244
rect 19616 4004 19668 4010
rect 19616 3946 19668 3952
rect 19340 3528 19392 3534
rect 19340 3470 19392 3476
rect 17592 3188 17644 3194
rect 17592 3130 17644 3136
rect 19628 2990 19656 3946
rect 19720 3466 19748 5238
rect 19996 5234 20024 8978
rect 20076 8900 20128 8906
rect 20076 8842 20128 8848
rect 20088 8362 20116 8842
rect 20628 8832 20680 8838
rect 20628 8774 20680 8780
rect 20640 8566 20668 8774
rect 20916 8634 20944 9522
rect 21468 9518 21496 10066
rect 21456 9512 21508 9518
rect 21456 9454 21508 9460
rect 21468 8974 21496 9454
rect 21456 8968 21508 8974
rect 21456 8910 21508 8916
rect 20904 8628 20956 8634
rect 20904 8570 20956 8576
rect 20628 8560 20680 8566
rect 20628 8502 20680 8508
rect 21744 8514 21772 10610
rect 21928 9926 21956 10950
rect 22296 10742 22324 11290
rect 22664 11218 22692 11562
rect 22652 11212 22704 11218
rect 22652 11154 22704 11160
rect 23388 11212 23440 11218
rect 23388 11154 23440 11160
rect 22560 10804 22612 10810
rect 22560 10746 22612 10752
rect 22284 10736 22336 10742
rect 22284 10678 22336 10684
rect 22572 10062 22600 10746
rect 22744 10736 22796 10742
rect 22744 10678 22796 10684
rect 22756 10266 22784 10678
rect 22744 10260 22796 10266
rect 22744 10202 22796 10208
rect 23400 10198 23428 11154
rect 23848 11076 23900 11082
rect 23848 11018 23900 11024
rect 23860 10470 23888 11018
rect 24214 10908 24522 10917
rect 24214 10906 24220 10908
rect 24276 10906 24300 10908
rect 24356 10906 24380 10908
rect 24436 10906 24460 10908
rect 24516 10906 24522 10908
rect 24276 10854 24278 10906
rect 24458 10854 24460 10906
rect 24214 10852 24220 10854
rect 24276 10852 24300 10854
rect 24356 10852 24380 10854
rect 24436 10852 24460 10854
rect 24516 10852 24522 10854
rect 24214 10843 24522 10852
rect 23848 10464 23900 10470
rect 23848 10406 23900 10412
rect 23388 10192 23440 10198
rect 23388 10134 23440 10140
rect 22560 10056 22612 10062
rect 22560 9998 22612 10004
rect 21916 9920 21968 9926
rect 21916 9862 21968 9868
rect 21824 8900 21876 8906
rect 21824 8842 21876 8848
rect 21836 8634 21864 8842
rect 21824 8628 21876 8634
rect 21824 8570 21876 8576
rect 21744 8498 21864 8514
rect 20812 8492 20864 8498
rect 21744 8492 21876 8498
rect 21744 8486 21824 8492
rect 20812 8434 20864 8440
rect 21824 8434 21876 8440
rect 20076 8356 20128 8362
rect 20076 8298 20128 8304
rect 20088 7410 20116 8298
rect 20720 8288 20772 8294
rect 20720 8230 20772 8236
rect 20214 8188 20522 8197
rect 20214 8186 20220 8188
rect 20276 8186 20300 8188
rect 20356 8186 20380 8188
rect 20436 8186 20460 8188
rect 20516 8186 20522 8188
rect 20276 8134 20278 8186
rect 20458 8134 20460 8186
rect 20214 8132 20220 8134
rect 20276 8132 20300 8134
rect 20356 8132 20380 8134
rect 20436 8132 20460 8134
rect 20516 8132 20522 8134
rect 20214 8123 20522 8132
rect 20352 7880 20404 7886
rect 20352 7822 20404 7828
rect 20364 7546 20392 7822
rect 20352 7540 20404 7546
rect 20352 7482 20404 7488
rect 20076 7404 20128 7410
rect 20076 7346 20128 7352
rect 20732 7342 20760 8230
rect 20824 7546 20852 8434
rect 20996 8288 21048 8294
rect 20996 8230 21048 8236
rect 21008 7954 21036 8230
rect 20996 7948 21048 7954
rect 20996 7890 21048 7896
rect 21088 7744 21140 7750
rect 21088 7686 21140 7692
rect 21100 7546 21128 7686
rect 20812 7540 20864 7546
rect 20812 7482 20864 7488
rect 21088 7540 21140 7546
rect 21088 7482 21140 7488
rect 20720 7336 20772 7342
rect 20720 7278 20772 7284
rect 20214 7100 20522 7109
rect 20214 7098 20220 7100
rect 20276 7098 20300 7100
rect 20356 7098 20380 7100
rect 20436 7098 20460 7100
rect 20516 7098 20522 7100
rect 20276 7046 20278 7098
rect 20458 7046 20460 7098
rect 20214 7044 20220 7046
rect 20276 7044 20300 7046
rect 20356 7044 20380 7046
rect 20436 7044 20460 7046
rect 20516 7044 20522 7046
rect 20214 7035 20522 7044
rect 21100 6458 21128 7482
rect 21836 7410 21864 8434
rect 21928 7546 21956 9862
rect 22572 9722 22600 9998
rect 22744 9920 22796 9926
rect 22744 9862 22796 9868
rect 22560 9716 22612 9722
rect 22560 9658 22612 9664
rect 22756 9586 22784 9862
rect 22100 9580 22152 9586
rect 22100 9522 22152 9528
rect 22744 9580 22796 9586
rect 22744 9522 22796 9528
rect 23020 9580 23072 9586
rect 23020 9522 23072 9528
rect 22112 9178 22140 9522
rect 23032 9466 23060 9522
rect 23032 9438 23152 9466
rect 22836 9376 22888 9382
rect 22836 9318 22888 9324
rect 22100 9172 22152 9178
rect 22100 9114 22152 9120
rect 22848 9042 22876 9318
rect 23124 9042 23152 9438
rect 23400 9042 23428 10134
rect 23480 9716 23532 9722
rect 23480 9658 23532 9664
rect 22836 9036 22888 9042
rect 22836 8978 22888 8984
rect 23112 9036 23164 9042
rect 23112 8978 23164 8984
rect 23388 9036 23440 9042
rect 23388 8978 23440 8984
rect 23124 8498 23152 8978
rect 23492 8906 23520 9658
rect 23480 8900 23532 8906
rect 23480 8842 23532 8848
rect 23112 8492 23164 8498
rect 23112 8434 23164 8440
rect 22008 8424 22060 8430
rect 22008 8366 22060 8372
rect 21916 7540 21968 7546
rect 21916 7482 21968 7488
rect 22020 7410 22048 8366
rect 22928 8288 22980 8294
rect 22928 8230 22980 8236
rect 22376 7948 22428 7954
rect 22376 7890 22428 7896
rect 22388 7410 22416 7890
rect 22560 7812 22612 7818
rect 22560 7754 22612 7760
rect 22572 7478 22600 7754
rect 22652 7744 22704 7750
rect 22652 7686 22704 7692
rect 22664 7478 22692 7686
rect 22940 7478 22968 8230
rect 23124 8022 23152 8434
rect 23492 8294 23520 8842
rect 23572 8560 23624 8566
rect 23572 8502 23624 8508
rect 23480 8288 23532 8294
rect 23480 8230 23532 8236
rect 23112 8016 23164 8022
rect 23112 7958 23164 7964
rect 23492 7886 23520 8230
rect 23584 8090 23612 8502
rect 23664 8424 23716 8430
rect 23664 8366 23716 8372
rect 23676 8090 23704 8366
rect 23572 8084 23624 8090
rect 23572 8026 23624 8032
rect 23664 8084 23716 8090
rect 23664 8026 23716 8032
rect 23112 7880 23164 7886
rect 23112 7822 23164 7828
rect 23480 7880 23532 7886
rect 23480 7822 23532 7828
rect 22560 7472 22612 7478
rect 22560 7414 22612 7420
rect 22652 7472 22704 7478
rect 22652 7414 22704 7420
rect 22928 7472 22980 7478
rect 22928 7414 22980 7420
rect 21824 7404 21876 7410
rect 21824 7346 21876 7352
rect 22008 7404 22060 7410
rect 22008 7346 22060 7352
rect 22376 7404 22428 7410
rect 22376 7346 22428 7352
rect 21916 7200 21968 7206
rect 21916 7142 21968 7148
rect 21364 6860 21416 6866
rect 21364 6802 21416 6808
rect 21376 6458 21404 6802
rect 21928 6730 21956 7142
rect 22388 7002 22416 7346
rect 22376 6996 22428 7002
rect 22376 6938 22428 6944
rect 21916 6724 21968 6730
rect 21916 6666 21968 6672
rect 22100 6656 22152 6662
rect 22100 6598 22152 6604
rect 21088 6452 21140 6458
rect 21088 6394 21140 6400
rect 21364 6452 21416 6458
rect 21364 6394 21416 6400
rect 22112 6322 22140 6598
rect 22388 6390 22416 6938
rect 22376 6384 22428 6390
rect 22376 6326 22428 6332
rect 22100 6316 22152 6322
rect 22100 6258 22152 6264
rect 20628 6248 20680 6254
rect 20628 6190 20680 6196
rect 20904 6248 20956 6254
rect 20904 6190 20956 6196
rect 22376 6248 22428 6254
rect 22376 6190 22428 6196
rect 20214 6012 20522 6021
rect 20214 6010 20220 6012
rect 20276 6010 20300 6012
rect 20356 6010 20380 6012
rect 20436 6010 20460 6012
rect 20516 6010 20522 6012
rect 20276 5958 20278 6010
rect 20458 5958 20460 6010
rect 20214 5956 20220 5958
rect 20276 5956 20300 5958
rect 20356 5956 20380 5958
rect 20436 5956 20460 5958
rect 20516 5956 20522 5958
rect 20214 5947 20522 5956
rect 20640 5574 20668 6190
rect 20812 5636 20864 5642
rect 20812 5578 20864 5584
rect 20168 5568 20220 5574
rect 20168 5510 20220 5516
rect 20628 5568 20680 5574
rect 20628 5510 20680 5516
rect 20180 5370 20208 5510
rect 20824 5370 20852 5578
rect 20168 5364 20220 5370
rect 20168 5306 20220 5312
rect 20812 5364 20864 5370
rect 20812 5306 20864 5312
rect 19984 5228 20036 5234
rect 19984 5170 20036 5176
rect 20628 5228 20680 5234
rect 20628 5170 20680 5176
rect 19800 4616 19852 4622
rect 19800 4558 19852 4564
rect 19812 3942 19840 4558
rect 19892 4480 19944 4486
rect 19892 4422 19944 4428
rect 19904 3942 19932 4422
rect 19800 3936 19852 3942
rect 19800 3878 19852 3884
rect 19892 3936 19944 3942
rect 19892 3878 19944 3884
rect 19708 3460 19760 3466
rect 19708 3402 19760 3408
rect 19720 3058 19748 3402
rect 19812 3058 19840 3878
rect 19708 3052 19760 3058
rect 19708 2994 19760 3000
rect 19800 3052 19852 3058
rect 19800 2994 19852 3000
rect 17224 2984 17276 2990
rect 17224 2926 17276 2932
rect 19616 2984 19668 2990
rect 19616 2926 19668 2932
rect 17040 2916 17092 2922
rect 17040 2858 17092 2864
rect 17236 2802 17264 2926
rect 18512 2916 18564 2922
rect 18512 2858 18564 2864
rect 16212 2644 16264 2650
rect 16212 2586 16264 2592
rect 15660 2508 15712 2514
rect 15660 2450 15712 2456
rect 15936 2508 15988 2514
rect 15936 2450 15988 2456
rect 16592 2446 16620 2790
rect 16960 2774 17264 2802
rect 18420 2848 18472 2854
rect 18420 2790 18472 2796
rect 16672 2508 16724 2514
rect 16672 2450 16724 2456
rect 16580 2440 16632 2446
rect 16580 2382 16632 2388
rect 16214 2204 16522 2213
rect 16214 2202 16220 2204
rect 16276 2202 16300 2204
rect 16356 2202 16380 2204
rect 16436 2202 16460 2204
rect 16516 2202 16522 2204
rect 16276 2150 16278 2202
rect 16458 2150 16460 2202
rect 16214 2148 16220 2150
rect 16276 2148 16300 2150
rect 16356 2148 16380 2150
rect 16436 2148 16460 2150
rect 16516 2148 16522 2150
rect 16214 2139 16522 2148
rect 16684 2106 16712 2450
rect 18432 2446 18460 2790
rect 18420 2440 18472 2446
rect 18420 2382 18472 2388
rect 17776 2372 17828 2378
rect 17776 2314 17828 2320
rect 17500 2304 17552 2310
rect 17500 2246 17552 2252
rect 16672 2100 16724 2106
rect 16672 2042 16724 2048
rect 17512 2038 17540 2246
rect 17788 2106 17816 2314
rect 18524 2106 18552 2858
rect 19628 2446 19656 2926
rect 19904 2514 19932 3878
rect 19996 2514 20024 5170
rect 20076 5160 20128 5166
rect 20076 5102 20128 5108
rect 20088 3924 20116 5102
rect 20214 4924 20522 4933
rect 20214 4922 20220 4924
rect 20276 4922 20300 4924
rect 20356 4922 20380 4924
rect 20436 4922 20460 4924
rect 20516 4922 20522 4924
rect 20276 4870 20278 4922
rect 20458 4870 20460 4922
rect 20214 4868 20220 4870
rect 20276 4868 20300 4870
rect 20356 4868 20380 4870
rect 20436 4868 20460 4870
rect 20516 4868 20522 4870
rect 20214 4859 20522 4868
rect 20352 4480 20404 4486
rect 20352 4422 20404 4428
rect 20364 4146 20392 4422
rect 20640 4282 20668 5170
rect 20720 5024 20772 5030
rect 20720 4966 20772 4972
rect 20732 4690 20760 4966
rect 20916 4826 20944 6190
rect 22388 5370 22416 6190
rect 22376 5364 22428 5370
rect 22376 5306 22428 5312
rect 22388 4826 22416 5306
rect 20904 4820 20956 4826
rect 20904 4762 20956 4768
rect 22376 4820 22428 4826
rect 22376 4762 22428 4768
rect 20720 4684 20772 4690
rect 20720 4626 20772 4632
rect 22572 4622 22600 7414
rect 23124 7002 23152 7822
rect 23112 6996 23164 7002
rect 23112 6938 23164 6944
rect 22652 6860 22704 6866
rect 22652 6802 22704 6808
rect 22664 6254 22692 6802
rect 23664 6384 23716 6390
rect 23664 6326 23716 6332
rect 23112 6316 23164 6322
rect 23112 6258 23164 6264
rect 22652 6248 22704 6254
rect 22652 6190 22704 6196
rect 22664 5166 22692 6190
rect 23124 5234 23152 6258
rect 23676 5914 23704 6326
rect 23664 5908 23716 5914
rect 23664 5850 23716 5856
rect 23388 5704 23440 5710
rect 23388 5646 23440 5652
rect 23572 5704 23624 5710
rect 23572 5646 23624 5652
rect 23756 5704 23808 5710
rect 23756 5646 23808 5652
rect 23296 5568 23348 5574
rect 23296 5510 23348 5516
rect 23112 5228 23164 5234
rect 23032 5188 23112 5216
rect 22652 5160 22704 5166
rect 22652 5102 22704 5108
rect 22560 4616 22612 4622
rect 22560 4558 22612 4564
rect 20996 4548 21048 4554
rect 20996 4490 21048 4496
rect 20628 4276 20680 4282
rect 20628 4218 20680 4224
rect 20352 4140 20404 4146
rect 20352 4082 20404 4088
rect 20364 3924 20392 4082
rect 20088 3896 20392 3924
rect 20088 3534 20116 3896
rect 20214 3836 20522 3845
rect 20214 3834 20220 3836
rect 20276 3834 20300 3836
rect 20356 3834 20380 3836
rect 20436 3834 20460 3836
rect 20516 3834 20522 3836
rect 20276 3782 20278 3834
rect 20458 3782 20460 3834
rect 20214 3780 20220 3782
rect 20276 3780 20300 3782
rect 20356 3780 20380 3782
rect 20436 3780 20460 3782
rect 20516 3780 20522 3782
rect 20214 3771 20522 3780
rect 20640 3738 20668 4218
rect 20812 4140 20864 4146
rect 20812 4082 20864 4088
rect 20628 3732 20680 3738
rect 20628 3674 20680 3680
rect 20824 3618 20852 4082
rect 21008 4010 21036 4490
rect 22560 4480 22612 4486
rect 22560 4422 22612 4428
rect 22572 4214 22600 4422
rect 22560 4208 22612 4214
rect 22560 4150 22612 4156
rect 23032 4146 23060 5188
rect 23112 5170 23164 5176
rect 23112 5092 23164 5098
rect 23112 5034 23164 5040
rect 23124 4826 23152 5034
rect 23112 4820 23164 4826
rect 23112 4762 23164 4768
rect 23020 4140 23072 4146
rect 23020 4082 23072 4088
rect 20996 4004 21048 4010
rect 20996 3946 21048 3952
rect 20640 3590 20852 3618
rect 21088 3664 21140 3670
rect 21088 3606 21140 3612
rect 20076 3528 20128 3534
rect 20076 3470 20128 3476
rect 20640 3466 20668 3590
rect 20628 3460 20680 3466
rect 20628 3402 20680 3408
rect 20076 2984 20128 2990
rect 20076 2926 20128 2932
rect 19892 2508 19944 2514
rect 19892 2450 19944 2456
rect 19984 2508 20036 2514
rect 19984 2450 20036 2456
rect 19616 2440 19668 2446
rect 19616 2382 19668 2388
rect 19064 2304 19116 2310
rect 19064 2246 19116 2252
rect 19708 2304 19760 2310
rect 19708 2246 19760 2252
rect 17776 2100 17828 2106
rect 17776 2042 17828 2048
rect 18512 2100 18564 2106
rect 18512 2042 18564 2048
rect 17500 2032 17552 2038
rect 17500 1974 17552 1980
rect 17788 1902 17816 2042
rect 17040 1896 17092 1902
rect 17040 1838 17092 1844
rect 17776 1896 17828 1902
rect 17776 1838 17828 1844
rect 17052 1562 17080 1838
rect 17040 1556 17092 1562
rect 17040 1498 17092 1504
rect 18524 1358 18552 2042
rect 19076 2038 19104 2246
rect 19064 2032 19116 2038
rect 19064 1974 19116 1980
rect 19720 1766 19748 2246
rect 19708 1760 19760 1766
rect 19708 1702 19760 1708
rect 19720 1426 19748 1702
rect 20088 1442 20116 2926
rect 20214 2748 20522 2757
rect 20214 2746 20220 2748
rect 20276 2746 20300 2748
rect 20356 2746 20380 2748
rect 20436 2746 20460 2748
rect 20516 2746 20522 2748
rect 20276 2694 20278 2746
rect 20458 2694 20460 2746
rect 20214 2692 20220 2694
rect 20276 2692 20300 2694
rect 20356 2692 20380 2694
rect 20436 2692 20460 2694
rect 20516 2692 20522 2694
rect 20214 2683 20522 2692
rect 20640 2446 20668 3402
rect 21100 3126 21128 3606
rect 23032 3602 23060 4082
rect 23308 4078 23336 5510
rect 23400 4826 23428 5646
rect 23388 4820 23440 4826
rect 23388 4762 23440 4768
rect 23296 4072 23348 4078
rect 23296 4014 23348 4020
rect 23020 3596 23072 3602
rect 23020 3538 23072 3544
rect 23584 3534 23612 5646
rect 23664 5296 23716 5302
rect 23664 5238 23716 5244
rect 23676 3738 23704 5238
rect 23768 4690 23796 5646
rect 23860 4690 23888 10406
rect 24124 10056 24176 10062
rect 24124 9998 24176 10004
rect 24136 8974 24164 9998
rect 24768 9988 24820 9994
rect 24768 9930 24820 9936
rect 24214 9820 24522 9829
rect 24214 9818 24220 9820
rect 24276 9818 24300 9820
rect 24356 9818 24380 9820
rect 24436 9818 24460 9820
rect 24516 9818 24522 9820
rect 24276 9766 24278 9818
rect 24458 9766 24460 9818
rect 24214 9764 24220 9766
rect 24276 9764 24300 9766
rect 24356 9764 24380 9766
rect 24436 9764 24460 9766
rect 24516 9764 24522 9766
rect 24214 9755 24522 9764
rect 24400 9580 24452 9586
rect 24400 9522 24452 9528
rect 24412 9178 24440 9522
rect 24780 9518 24808 9930
rect 24768 9512 24820 9518
rect 24768 9454 24820 9460
rect 24400 9172 24452 9178
rect 24400 9114 24452 9120
rect 24124 8968 24176 8974
rect 24124 8910 24176 8916
rect 24124 8832 24176 8838
rect 24124 8774 24176 8780
rect 24032 8084 24084 8090
rect 24032 8026 24084 8032
rect 24044 7342 24072 8026
rect 24136 7546 24164 8774
rect 24214 8732 24522 8741
rect 24214 8730 24220 8732
rect 24276 8730 24300 8732
rect 24356 8730 24380 8732
rect 24436 8730 24460 8732
rect 24516 8730 24522 8732
rect 24276 8678 24278 8730
rect 24458 8678 24460 8730
rect 24214 8676 24220 8678
rect 24276 8676 24300 8678
rect 24356 8676 24380 8678
rect 24436 8676 24460 8678
rect 24516 8676 24522 8678
rect 24214 8667 24522 8676
rect 24780 7954 24808 9454
rect 25136 8288 25188 8294
rect 25136 8230 25188 8236
rect 24768 7948 24820 7954
rect 24768 7890 24820 7896
rect 25148 7886 25176 8230
rect 25136 7880 25188 7886
rect 25136 7822 25188 7828
rect 24214 7644 24522 7653
rect 24214 7642 24220 7644
rect 24276 7642 24300 7644
rect 24356 7642 24380 7644
rect 24436 7642 24460 7644
rect 24516 7642 24522 7644
rect 24276 7590 24278 7642
rect 24458 7590 24460 7642
rect 24214 7588 24220 7590
rect 24276 7588 24300 7590
rect 24356 7588 24380 7590
rect 24436 7588 24460 7590
rect 24516 7588 24522 7590
rect 24214 7579 24522 7588
rect 24124 7540 24176 7546
rect 24124 7482 24176 7488
rect 24032 7336 24084 7342
rect 24032 7278 24084 7284
rect 23940 7268 23992 7274
rect 23940 7210 23992 7216
rect 23952 6254 23980 7210
rect 23940 6248 23992 6254
rect 23940 6190 23992 6196
rect 24044 4690 24072 7278
rect 24136 6798 24164 7482
rect 24584 7404 24636 7410
rect 24584 7346 24636 7352
rect 24596 7002 24624 7346
rect 24584 6996 24636 7002
rect 24584 6938 24636 6944
rect 24952 6860 25004 6866
rect 24952 6802 25004 6808
rect 24124 6792 24176 6798
rect 24964 6746 24992 6802
rect 25148 6798 25176 7822
rect 24124 6734 24176 6740
rect 24872 6718 24992 6746
rect 25136 6792 25188 6798
rect 25136 6734 25188 6740
rect 24214 6556 24522 6565
rect 24214 6554 24220 6556
rect 24276 6554 24300 6556
rect 24356 6554 24380 6556
rect 24436 6554 24460 6556
rect 24516 6554 24522 6556
rect 24276 6502 24278 6554
rect 24458 6502 24460 6554
rect 24214 6500 24220 6502
rect 24276 6500 24300 6502
rect 24356 6500 24380 6502
rect 24436 6500 24460 6502
rect 24516 6500 24522 6502
rect 24214 6491 24522 6500
rect 24214 5468 24522 5477
rect 24214 5466 24220 5468
rect 24276 5466 24300 5468
rect 24356 5466 24380 5468
rect 24436 5466 24460 5468
rect 24516 5466 24522 5468
rect 24276 5414 24278 5466
rect 24458 5414 24460 5466
rect 24214 5412 24220 5414
rect 24276 5412 24300 5414
rect 24356 5412 24380 5414
rect 24436 5412 24460 5414
rect 24516 5412 24522 5414
rect 24214 5403 24522 5412
rect 24872 4826 24900 6718
rect 25044 6656 25096 6662
rect 25044 6598 25096 6604
rect 25056 6458 25084 6598
rect 25044 6452 25096 6458
rect 25044 6394 25096 6400
rect 26160 5545 26188 16458
rect 26424 16040 26476 16046
rect 26424 15982 26476 15988
rect 26146 5536 26202 5545
rect 26146 5471 26202 5480
rect 24952 5024 25004 5030
rect 24952 4966 25004 4972
rect 24860 4820 24912 4826
rect 24860 4762 24912 4768
rect 24964 4690 24992 4966
rect 23756 4684 23808 4690
rect 23756 4626 23808 4632
rect 23848 4684 23900 4690
rect 23848 4626 23900 4632
rect 24032 4684 24084 4690
rect 24032 4626 24084 4632
rect 24952 4684 25004 4690
rect 24952 4626 25004 4632
rect 23664 3732 23716 3738
rect 23664 3674 23716 3680
rect 23768 3534 23796 4626
rect 24768 4480 24820 4486
rect 24768 4422 24820 4428
rect 24214 4380 24522 4389
rect 24214 4378 24220 4380
rect 24276 4378 24300 4380
rect 24356 4378 24380 4380
rect 24436 4378 24460 4380
rect 24516 4378 24522 4380
rect 24276 4326 24278 4378
rect 24458 4326 24460 4378
rect 24214 4324 24220 4326
rect 24276 4324 24300 4326
rect 24356 4324 24380 4326
rect 24436 4324 24460 4326
rect 24516 4324 24522 4326
rect 24214 4315 24522 4324
rect 24780 4282 24808 4422
rect 24768 4276 24820 4282
rect 24768 4218 24820 4224
rect 23572 3528 23624 3534
rect 23572 3470 23624 3476
rect 23756 3528 23808 3534
rect 23756 3470 23808 3476
rect 22008 3460 22060 3466
rect 22008 3402 22060 3408
rect 21456 3392 21508 3398
rect 21456 3334 21508 3340
rect 21548 3392 21600 3398
rect 21548 3334 21600 3340
rect 21088 3120 21140 3126
rect 21088 3062 21140 3068
rect 21468 3058 21496 3334
rect 21560 3194 21588 3334
rect 22020 3194 22048 3402
rect 21548 3188 21600 3194
rect 21548 3130 21600 3136
rect 22008 3188 22060 3194
rect 22008 3130 22060 3136
rect 23768 3058 23796 3470
rect 24214 3292 24522 3301
rect 24214 3290 24220 3292
rect 24276 3290 24300 3292
rect 24356 3290 24380 3292
rect 24436 3290 24460 3292
rect 24516 3290 24522 3292
rect 24276 3238 24278 3290
rect 24458 3238 24460 3290
rect 24214 3236 24220 3238
rect 24276 3236 24300 3238
rect 24356 3236 24380 3238
rect 24436 3236 24460 3238
rect 24516 3236 24522 3238
rect 24214 3227 24522 3236
rect 21456 3052 21508 3058
rect 21456 2994 21508 3000
rect 23756 3052 23808 3058
rect 23756 2994 23808 3000
rect 20628 2440 20680 2446
rect 20628 2382 20680 2388
rect 20444 2304 20496 2310
rect 20444 2246 20496 2252
rect 20456 2038 20484 2246
rect 24214 2204 24522 2213
rect 24214 2202 24220 2204
rect 24276 2202 24300 2204
rect 24356 2202 24380 2204
rect 24436 2202 24460 2204
rect 24516 2202 24522 2204
rect 24276 2150 24278 2202
rect 24458 2150 24460 2202
rect 24214 2148 24220 2150
rect 24276 2148 24300 2150
rect 24356 2148 24380 2150
rect 24436 2148 24460 2150
rect 24516 2148 24522 2150
rect 24214 2139 24522 2148
rect 20444 2032 20496 2038
rect 20444 1974 20496 1980
rect 26146 2000 26202 2009
rect 26436 1986 26464 15982
rect 26202 1958 26464 1986
rect 26146 1935 26202 1944
rect 20214 1660 20522 1669
rect 20214 1658 20220 1660
rect 20276 1658 20300 1660
rect 20356 1658 20380 1660
rect 20436 1658 20460 1660
rect 20516 1658 20522 1660
rect 20276 1606 20278 1658
rect 20458 1606 20460 1658
rect 20214 1604 20220 1606
rect 20276 1604 20300 1606
rect 20356 1604 20380 1606
rect 20436 1604 20460 1606
rect 20516 1604 20522 1606
rect 20214 1595 20522 1604
rect 19708 1420 19760 1426
rect 20088 1414 20208 1442
rect 19708 1362 19760 1368
rect 18512 1352 18564 1358
rect 18512 1294 18564 1300
rect 15108 1284 15160 1290
rect 15108 1226 15160 1232
rect 14556 1216 14608 1222
rect 6656 1142 6776 1170
rect 14556 1158 14608 1164
rect 6748 800 6776 1142
rect 8214 1116 8522 1125
rect 8214 1114 8220 1116
rect 8276 1114 8300 1116
rect 8356 1114 8380 1116
rect 8436 1114 8460 1116
rect 8516 1114 8522 1116
rect 8276 1062 8278 1114
rect 8458 1062 8460 1114
rect 8214 1060 8220 1062
rect 8276 1060 8300 1062
rect 8356 1060 8380 1062
rect 8436 1060 8460 1062
rect 8516 1060 8522 1062
rect 8214 1051 8522 1060
rect 16214 1116 16522 1125
rect 16214 1114 16220 1116
rect 16276 1114 16300 1116
rect 16356 1114 16380 1116
rect 16436 1114 16460 1116
rect 16516 1114 16522 1116
rect 16276 1062 16278 1114
rect 16458 1062 16460 1114
rect 16214 1060 16220 1062
rect 16276 1060 16300 1062
rect 16356 1060 16380 1062
rect 16436 1060 16460 1062
rect 16516 1060 16522 1062
rect 16214 1051 16522 1060
rect 20180 800 20208 1414
rect 24214 1116 24522 1125
rect 24214 1114 24220 1116
rect 24276 1114 24300 1116
rect 24356 1114 24380 1116
rect 24436 1114 24460 1116
rect 24516 1114 24522 1116
rect 24276 1062 24278 1114
rect 24458 1062 24460 1114
rect 24214 1060 24220 1062
rect 24276 1060 24300 1062
rect 24356 1060 24380 1062
rect 24436 1060 24460 1062
rect 24516 1060 24522 1062
rect 24214 1051 24522 1060
rect 6734 0 6790 800
rect 20166 0 20222 800
<< via2 >>
rect 6734 20712 6790 20768
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4618 19624 4674 19680
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 3974 18536 4030 18592
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 5630 17448 5686 17504
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 8220 20698 8276 20700
rect 8300 20698 8356 20700
rect 8380 20698 8436 20700
rect 8460 20698 8516 20700
rect 8220 20646 8266 20698
rect 8266 20646 8276 20698
rect 8300 20646 8330 20698
rect 8330 20646 8342 20698
rect 8342 20646 8356 20698
rect 8380 20646 8394 20698
rect 8394 20646 8406 20698
rect 8406 20646 8436 20698
rect 8460 20646 8470 20698
rect 8470 20646 8516 20698
rect 8220 20644 8276 20646
rect 8300 20644 8356 20646
rect 8380 20644 8436 20646
rect 8460 20644 8516 20646
rect 8220 19610 8276 19612
rect 8300 19610 8356 19612
rect 8380 19610 8436 19612
rect 8460 19610 8516 19612
rect 8220 19558 8266 19610
rect 8266 19558 8276 19610
rect 8300 19558 8330 19610
rect 8330 19558 8342 19610
rect 8342 19558 8356 19610
rect 8380 19558 8394 19610
rect 8394 19558 8406 19610
rect 8406 19558 8436 19610
rect 8460 19558 8470 19610
rect 8470 19558 8516 19610
rect 8220 19556 8276 19558
rect 8300 19556 8356 19558
rect 8380 19556 8436 19558
rect 8460 19556 8516 19558
rect 7378 16360 7434 16416
rect 8220 18522 8276 18524
rect 8300 18522 8356 18524
rect 8380 18522 8436 18524
rect 8460 18522 8516 18524
rect 8220 18470 8266 18522
rect 8266 18470 8276 18522
rect 8300 18470 8330 18522
rect 8330 18470 8342 18522
rect 8342 18470 8356 18522
rect 8380 18470 8394 18522
rect 8394 18470 8406 18522
rect 8406 18470 8436 18522
rect 8460 18470 8470 18522
rect 8470 18470 8516 18522
rect 8220 18468 8276 18470
rect 8300 18468 8356 18470
rect 8380 18468 8436 18470
rect 8460 18468 8516 18470
rect 8220 17434 8276 17436
rect 8300 17434 8356 17436
rect 8380 17434 8436 17436
rect 8460 17434 8516 17436
rect 8220 17382 8266 17434
rect 8266 17382 8276 17434
rect 8300 17382 8330 17434
rect 8330 17382 8342 17434
rect 8342 17382 8356 17434
rect 8380 17382 8394 17434
rect 8394 17382 8406 17434
rect 8406 17382 8436 17434
rect 8460 17382 8470 17434
rect 8470 17382 8516 17434
rect 8220 17380 8276 17382
rect 8300 17380 8356 17382
rect 8380 17380 8436 17382
rect 8460 17380 8516 17382
rect 6918 15272 6974 15328
rect 6458 14184 6514 14240
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 1306 10920 1362 10976
rect 1306 8744 1362 8800
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 9218 17312 9274 17368
rect 8220 16346 8276 16348
rect 8300 16346 8356 16348
rect 8380 16346 8436 16348
rect 8460 16346 8516 16348
rect 8220 16294 8266 16346
rect 8266 16294 8276 16346
rect 8300 16294 8330 16346
rect 8330 16294 8342 16346
rect 8342 16294 8356 16346
rect 8380 16294 8394 16346
rect 8394 16294 8406 16346
rect 8406 16294 8436 16346
rect 8460 16294 8470 16346
rect 8470 16294 8516 16346
rect 8220 16292 8276 16294
rect 8300 16292 8356 16294
rect 8380 16292 8436 16294
rect 8460 16292 8516 16294
rect 10782 19760 10838 19816
rect 12220 20154 12276 20156
rect 12300 20154 12356 20156
rect 12380 20154 12436 20156
rect 12460 20154 12516 20156
rect 12220 20102 12266 20154
rect 12266 20102 12276 20154
rect 12300 20102 12330 20154
rect 12330 20102 12342 20154
rect 12342 20102 12356 20154
rect 12380 20102 12394 20154
rect 12394 20102 12406 20154
rect 12406 20102 12436 20154
rect 12460 20102 12470 20154
rect 12470 20102 12516 20154
rect 12220 20100 12276 20102
rect 12300 20100 12356 20102
rect 12380 20100 12436 20102
rect 12460 20100 12516 20102
rect 8220 15258 8276 15260
rect 8300 15258 8356 15260
rect 8380 15258 8436 15260
rect 8460 15258 8516 15260
rect 8220 15206 8266 15258
rect 8266 15206 8276 15258
rect 8300 15206 8330 15258
rect 8330 15206 8342 15258
rect 8342 15206 8356 15258
rect 8380 15206 8394 15258
rect 8394 15206 8406 15258
rect 8406 15206 8436 15258
rect 8460 15206 8470 15258
rect 8470 15206 8516 15258
rect 8220 15204 8276 15206
rect 8300 15204 8356 15206
rect 8380 15204 8436 15206
rect 8460 15204 8516 15206
rect 8220 14170 8276 14172
rect 8300 14170 8356 14172
rect 8380 14170 8436 14172
rect 8460 14170 8516 14172
rect 8220 14118 8266 14170
rect 8266 14118 8276 14170
rect 8300 14118 8330 14170
rect 8330 14118 8342 14170
rect 8342 14118 8356 14170
rect 8380 14118 8394 14170
rect 8394 14118 8406 14170
rect 8406 14118 8436 14170
rect 8460 14118 8470 14170
rect 8470 14118 8516 14170
rect 8220 14116 8276 14118
rect 8300 14116 8356 14118
rect 8380 14116 8436 14118
rect 8460 14116 8516 14118
rect 10414 18128 10470 18184
rect 10138 17448 10194 17504
rect 9862 17040 9918 17096
rect 10230 17176 10286 17232
rect 9770 16360 9826 16416
rect 8220 13082 8276 13084
rect 8300 13082 8356 13084
rect 8380 13082 8436 13084
rect 8460 13082 8516 13084
rect 8220 13030 8266 13082
rect 8266 13030 8276 13082
rect 8300 13030 8330 13082
rect 8330 13030 8342 13082
rect 8342 13030 8356 13082
rect 8380 13030 8394 13082
rect 8394 13030 8406 13082
rect 8406 13030 8436 13082
rect 8460 13030 8470 13082
rect 8470 13030 8516 13082
rect 8220 13028 8276 13030
rect 8300 13028 8356 13030
rect 8380 13028 8436 13030
rect 8460 13028 8516 13030
rect 10966 18264 11022 18320
rect 10874 17720 10930 17776
rect 10690 17584 10746 17640
rect 10598 17196 10654 17232
rect 10598 17176 10600 17196
rect 10600 17176 10652 17196
rect 10652 17176 10654 17196
rect 10414 16632 10470 16688
rect 6182 9832 6238 9888
rect 3330 6568 3386 6624
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 3054 5480 3110 5536
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4986 7656 5042 7712
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 202 2488 258 2544
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 5078 4392 5134 4448
rect 4220 1658 4276 1660
rect 4300 1658 4356 1660
rect 4380 1658 4436 1660
rect 4460 1658 4516 1660
rect 4220 1606 4266 1658
rect 4266 1606 4276 1658
rect 4300 1606 4330 1658
rect 4330 1606 4342 1658
rect 4342 1606 4356 1658
rect 4380 1606 4394 1658
rect 4394 1606 4406 1658
rect 4406 1606 4436 1658
rect 4460 1606 4470 1658
rect 4470 1606 4516 1658
rect 4220 1604 4276 1606
rect 4300 1604 4356 1606
rect 4380 1604 4436 1606
rect 4460 1604 4516 1606
rect 8220 11994 8276 11996
rect 8300 11994 8356 11996
rect 8380 11994 8436 11996
rect 8460 11994 8516 11996
rect 8220 11942 8266 11994
rect 8266 11942 8276 11994
rect 8300 11942 8330 11994
rect 8330 11942 8342 11994
rect 8342 11942 8356 11994
rect 8380 11942 8394 11994
rect 8394 11942 8406 11994
rect 8406 11942 8436 11994
rect 8460 11942 8470 11994
rect 8470 11942 8516 11994
rect 8220 11940 8276 11942
rect 8300 11940 8356 11942
rect 8380 11940 8436 11942
rect 8460 11940 8516 11942
rect 10966 16088 11022 16144
rect 11610 19080 11666 19136
rect 11702 18808 11758 18864
rect 11334 18672 11390 18728
rect 11426 18536 11482 18592
rect 11426 18400 11482 18456
rect 11610 17856 11666 17912
rect 11242 16496 11298 16552
rect 11794 17484 11796 17504
rect 11796 17484 11848 17504
rect 11848 17484 11850 17504
rect 11794 17448 11850 17484
rect 12220 19066 12276 19068
rect 12300 19066 12356 19068
rect 12380 19066 12436 19068
rect 12460 19066 12516 19068
rect 12220 19014 12266 19066
rect 12266 19014 12276 19066
rect 12300 19014 12330 19066
rect 12330 19014 12342 19066
rect 12342 19014 12356 19066
rect 12380 19014 12394 19066
rect 12394 19014 12406 19066
rect 12406 19014 12436 19066
rect 12460 19014 12470 19066
rect 12470 19014 12516 19066
rect 12220 19012 12276 19014
rect 12300 19012 12356 19014
rect 12380 19012 12436 19014
rect 12460 19012 12516 19014
rect 12070 18844 12072 18864
rect 12072 18844 12124 18864
rect 12124 18844 12126 18864
rect 12070 18808 12126 18844
rect 12438 18808 12494 18864
rect 12622 18708 12624 18728
rect 12624 18708 12676 18728
rect 12676 18708 12678 18728
rect 12622 18672 12678 18708
rect 12346 18420 12402 18456
rect 12346 18400 12348 18420
rect 12348 18400 12400 18420
rect 12400 18400 12402 18420
rect 12714 18284 12770 18320
rect 12714 18264 12716 18284
rect 12716 18264 12768 18284
rect 12768 18264 12770 18284
rect 12070 18128 12126 18184
rect 12220 17978 12276 17980
rect 12300 17978 12356 17980
rect 12380 17978 12436 17980
rect 12460 17978 12516 17980
rect 12220 17926 12266 17978
rect 12266 17926 12276 17978
rect 12300 17926 12330 17978
rect 12330 17926 12342 17978
rect 12342 17926 12356 17978
rect 12380 17926 12394 17978
rect 12394 17926 12406 17978
rect 12406 17926 12436 17978
rect 12460 17926 12470 17978
rect 12470 17926 12516 17978
rect 12220 17924 12276 17926
rect 12300 17924 12356 17926
rect 12380 17924 12436 17926
rect 12460 17924 12516 17926
rect 12898 17720 12954 17776
rect 13818 18808 13874 18864
rect 13450 18264 13506 18320
rect 12714 17312 12770 17368
rect 11610 16788 11666 16824
rect 11610 16768 11612 16788
rect 11612 16768 11664 16788
rect 11664 16768 11666 16788
rect 12070 16904 12126 16960
rect 12220 16890 12276 16892
rect 12300 16890 12356 16892
rect 12380 16890 12436 16892
rect 12460 16890 12516 16892
rect 12220 16838 12266 16890
rect 12266 16838 12276 16890
rect 12300 16838 12330 16890
rect 12330 16838 12342 16890
rect 12342 16838 12356 16890
rect 12380 16838 12394 16890
rect 12394 16838 12406 16890
rect 12406 16838 12436 16890
rect 12460 16838 12470 16890
rect 12470 16838 12516 16890
rect 12220 16836 12276 16838
rect 12300 16836 12356 16838
rect 12380 16836 12436 16838
rect 12460 16836 12516 16838
rect 12070 16632 12126 16688
rect 12162 16532 12164 16552
rect 12164 16532 12216 16552
rect 12216 16532 12218 16552
rect 12162 16496 12218 16532
rect 11610 16244 11666 16280
rect 11886 16360 11942 16416
rect 11610 16224 11612 16244
rect 11612 16224 11664 16244
rect 11664 16224 11666 16244
rect 12220 15802 12276 15804
rect 12300 15802 12356 15804
rect 12380 15802 12436 15804
rect 12460 15802 12516 15804
rect 12220 15750 12266 15802
rect 12266 15750 12276 15802
rect 12300 15750 12330 15802
rect 12330 15750 12342 15802
rect 12342 15750 12356 15802
rect 12380 15750 12394 15802
rect 12394 15750 12406 15802
rect 12406 15750 12436 15802
rect 12460 15750 12470 15802
rect 12470 15750 12516 15802
rect 12220 15748 12276 15750
rect 12300 15748 12356 15750
rect 12380 15748 12436 15750
rect 12460 15748 12516 15750
rect 13818 17604 13874 17640
rect 13818 17584 13820 17604
rect 13820 17584 13872 17604
rect 13872 17584 13874 17604
rect 13634 17448 13690 17504
rect 15474 18536 15530 18592
rect 16220 20698 16276 20700
rect 16300 20698 16356 20700
rect 16380 20698 16436 20700
rect 16460 20698 16516 20700
rect 16220 20646 16266 20698
rect 16266 20646 16276 20698
rect 16300 20646 16330 20698
rect 16330 20646 16342 20698
rect 16342 20646 16356 20698
rect 16380 20646 16394 20698
rect 16394 20646 16406 20698
rect 16406 20646 16436 20698
rect 16460 20646 16470 20698
rect 16470 20646 16516 20698
rect 16220 20644 16276 20646
rect 16300 20644 16356 20646
rect 16380 20644 16436 20646
rect 16460 20644 16516 20646
rect 16670 19760 16726 19816
rect 16220 19610 16276 19612
rect 16300 19610 16356 19612
rect 16380 19610 16436 19612
rect 16460 19610 16516 19612
rect 16220 19558 16266 19610
rect 16266 19558 16276 19610
rect 16300 19558 16330 19610
rect 16330 19558 16342 19610
rect 16342 19558 16356 19610
rect 16380 19558 16394 19610
rect 16394 19558 16406 19610
rect 16406 19558 16436 19610
rect 16460 19558 16470 19610
rect 16470 19558 16516 19610
rect 16220 19556 16276 19558
rect 16300 19556 16356 19558
rect 16380 19556 16436 19558
rect 16460 19556 16516 19558
rect 16220 18522 16276 18524
rect 16300 18522 16356 18524
rect 16380 18522 16436 18524
rect 16460 18522 16516 18524
rect 16220 18470 16266 18522
rect 16266 18470 16276 18522
rect 16300 18470 16330 18522
rect 16330 18470 16342 18522
rect 16342 18470 16356 18522
rect 16380 18470 16394 18522
rect 16394 18470 16406 18522
rect 16406 18470 16436 18522
rect 16460 18470 16470 18522
rect 16470 18470 16516 18522
rect 16220 18468 16276 18470
rect 16300 18468 16356 18470
rect 16380 18468 16436 18470
rect 16460 18468 16516 18470
rect 13542 17040 13598 17096
rect 15382 17176 15438 17232
rect 14462 16632 14518 16688
rect 5906 3304 5962 3360
rect 8220 10906 8276 10908
rect 8300 10906 8356 10908
rect 8380 10906 8436 10908
rect 8460 10906 8516 10908
rect 8220 10854 8266 10906
rect 8266 10854 8276 10906
rect 8300 10854 8330 10906
rect 8330 10854 8342 10906
rect 8342 10854 8356 10906
rect 8380 10854 8394 10906
rect 8394 10854 8406 10906
rect 8406 10854 8436 10906
rect 8460 10854 8470 10906
rect 8470 10854 8516 10906
rect 8220 10852 8276 10854
rect 8300 10852 8356 10854
rect 8380 10852 8436 10854
rect 8460 10852 8516 10854
rect 8220 9818 8276 9820
rect 8300 9818 8356 9820
rect 8380 9818 8436 9820
rect 8460 9818 8516 9820
rect 8220 9766 8266 9818
rect 8266 9766 8276 9818
rect 8300 9766 8330 9818
rect 8330 9766 8342 9818
rect 8342 9766 8356 9818
rect 8380 9766 8394 9818
rect 8394 9766 8406 9818
rect 8406 9766 8436 9818
rect 8460 9766 8470 9818
rect 8470 9766 8516 9818
rect 8220 9764 8276 9766
rect 8300 9764 8356 9766
rect 8380 9764 8436 9766
rect 8460 9764 8516 9766
rect 8220 8730 8276 8732
rect 8300 8730 8356 8732
rect 8380 8730 8436 8732
rect 8460 8730 8516 8732
rect 8220 8678 8266 8730
rect 8266 8678 8276 8730
rect 8300 8678 8330 8730
rect 8330 8678 8342 8730
rect 8342 8678 8356 8730
rect 8380 8678 8394 8730
rect 8394 8678 8406 8730
rect 8406 8678 8436 8730
rect 8460 8678 8470 8730
rect 8470 8678 8516 8730
rect 8220 8676 8276 8678
rect 8300 8676 8356 8678
rect 8380 8676 8436 8678
rect 8460 8676 8516 8678
rect 8220 7642 8276 7644
rect 8300 7642 8356 7644
rect 8380 7642 8436 7644
rect 8460 7642 8516 7644
rect 8220 7590 8266 7642
rect 8266 7590 8276 7642
rect 8300 7590 8330 7642
rect 8330 7590 8342 7642
rect 8342 7590 8356 7642
rect 8380 7590 8394 7642
rect 8394 7590 8406 7642
rect 8406 7590 8436 7642
rect 8460 7590 8470 7642
rect 8470 7590 8516 7642
rect 8220 7588 8276 7590
rect 8300 7588 8356 7590
rect 8380 7588 8436 7590
rect 8460 7588 8516 7590
rect 8220 6554 8276 6556
rect 8300 6554 8356 6556
rect 8380 6554 8436 6556
rect 8460 6554 8516 6556
rect 8220 6502 8266 6554
rect 8266 6502 8276 6554
rect 8300 6502 8330 6554
rect 8330 6502 8342 6554
rect 8342 6502 8356 6554
rect 8380 6502 8394 6554
rect 8394 6502 8406 6554
rect 8406 6502 8436 6554
rect 8460 6502 8470 6554
rect 8470 6502 8516 6554
rect 8220 6500 8276 6502
rect 8300 6500 8356 6502
rect 8380 6500 8436 6502
rect 8460 6500 8516 6502
rect 8220 5466 8276 5468
rect 8300 5466 8356 5468
rect 8380 5466 8436 5468
rect 8460 5466 8516 5468
rect 8220 5414 8266 5466
rect 8266 5414 8276 5466
rect 8300 5414 8330 5466
rect 8330 5414 8342 5466
rect 8342 5414 8356 5466
rect 8380 5414 8394 5466
rect 8394 5414 8406 5466
rect 8406 5414 8436 5466
rect 8460 5414 8470 5466
rect 8470 5414 8516 5466
rect 8220 5412 8276 5414
rect 8300 5412 8356 5414
rect 8380 5412 8436 5414
rect 8460 5412 8516 5414
rect 846 1264 902 1320
rect 8220 4378 8276 4380
rect 8300 4378 8356 4380
rect 8380 4378 8436 4380
rect 8460 4378 8516 4380
rect 8220 4326 8266 4378
rect 8266 4326 8276 4378
rect 8300 4326 8330 4378
rect 8330 4326 8342 4378
rect 8342 4326 8356 4378
rect 8380 4326 8394 4378
rect 8394 4326 8406 4378
rect 8406 4326 8436 4378
rect 8460 4326 8470 4378
rect 8470 4326 8516 4378
rect 8220 4324 8276 4326
rect 8300 4324 8356 4326
rect 8380 4324 8436 4326
rect 8460 4324 8516 4326
rect 8220 3290 8276 3292
rect 8300 3290 8356 3292
rect 8380 3290 8436 3292
rect 8460 3290 8516 3292
rect 8220 3238 8266 3290
rect 8266 3238 8276 3290
rect 8300 3238 8330 3290
rect 8330 3238 8342 3290
rect 8342 3238 8356 3290
rect 8380 3238 8394 3290
rect 8394 3238 8406 3290
rect 8406 3238 8436 3290
rect 8460 3238 8470 3290
rect 8470 3238 8516 3290
rect 8220 3236 8276 3238
rect 8300 3236 8356 3238
rect 8380 3236 8436 3238
rect 8460 3236 8516 3238
rect 12220 14714 12276 14716
rect 12300 14714 12356 14716
rect 12380 14714 12436 14716
rect 12460 14714 12516 14716
rect 12220 14662 12266 14714
rect 12266 14662 12276 14714
rect 12300 14662 12330 14714
rect 12330 14662 12342 14714
rect 12342 14662 12356 14714
rect 12380 14662 12394 14714
rect 12394 14662 12406 14714
rect 12406 14662 12436 14714
rect 12460 14662 12470 14714
rect 12470 14662 12516 14714
rect 12220 14660 12276 14662
rect 12300 14660 12356 14662
rect 12380 14660 12436 14662
rect 12460 14660 12516 14662
rect 12220 13626 12276 13628
rect 12300 13626 12356 13628
rect 12380 13626 12436 13628
rect 12460 13626 12516 13628
rect 12220 13574 12266 13626
rect 12266 13574 12276 13626
rect 12300 13574 12330 13626
rect 12330 13574 12342 13626
rect 12342 13574 12356 13626
rect 12380 13574 12394 13626
rect 12394 13574 12406 13626
rect 12406 13574 12436 13626
rect 12460 13574 12470 13626
rect 12470 13574 12516 13626
rect 12220 13572 12276 13574
rect 12300 13572 12356 13574
rect 12380 13572 12436 13574
rect 12460 13572 12516 13574
rect 13634 12824 13690 12880
rect 12220 12538 12276 12540
rect 12300 12538 12356 12540
rect 12380 12538 12436 12540
rect 12460 12538 12516 12540
rect 12220 12486 12266 12538
rect 12266 12486 12276 12538
rect 12300 12486 12330 12538
rect 12330 12486 12342 12538
rect 12342 12486 12356 12538
rect 12380 12486 12394 12538
rect 12394 12486 12406 12538
rect 12406 12486 12436 12538
rect 12460 12486 12470 12538
rect 12470 12486 12516 12538
rect 12220 12484 12276 12486
rect 12300 12484 12356 12486
rect 12380 12484 12436 12486
rect 12460 12484 12516 12486
rect 10690 12144 10746 12200
rect 8220 2202 8276 2204
rect 8300 2202 8356 2204
rect 8380 2202 8436 2204
rect 8460 2202 8516 2204
rect 8220 2150 8266 2202
rect 8266 2150 8276 2202
rect 8300 2150 8330 2202
rect 8330 2150 8342 2202
rect 8342 2150 8356 2202
rect 8380 2150 8394 2202
rect 8394 2150 8406 2202
rect 8406 2150 8436 2202
rect 8460 2150 8470 2202
rect 8470 2150 8516 2202
rect 8220 2148 8276 2150
rect 8300 2148 8356 2150
rect 8380 2148 8436 2150
rect 8460 2148 8516 2150
rect 12220 11450 12276 11452
rect 12300 11450 12356 11452
rect 12380 11450 12436 11452
rect 12460 11450 12516 11452
rect 12220 11398 12266 11450
rect 12266 11398 12276 11450
rect 12300 11398 12330 11450
rect 12330 11398 12342 11450
rect 12342 11398 12356 11450
rect 12380 11398 12394 11450
rect 12394 11398 12406 11450
rect 12406 11398 12436 11450
rect 12460 11398 12470 11450
rect 12470 11398 12516 11450
rect 12220 11396 12276 11398
rect 12300 11396 12356 11398
rect 12380 11396 12436 11398
rect 12460 11396 12516 11398
rect 12220 10362 12276 10364
rect 12300 10362 12356 10364
rect 12380 10362 12436 10364
rect 12460 10362 12516 10364
rect 12220 10310 12266 10362
rect 12266 10310 12276 10362
rect 12300 10310 12330 10362
rect 12330 10310 12342 10362
rect 12342 10310 12356 10362
rect 12380 10310 12394 10362
rect 12394 10310 12406 10362
rect 12406 10310 12436 10362
rect 12460 10310 12470 10362
rect 12470 10310 12516 10362
rect 12220 10308 12276 10310
rect 12300 10308 12356 10310
rect 12380 10308 12436 10310
rect 12460 10308 12516 10310
rect 12220 9274 12276 9276
rect 12300 9274 12356 9276
rect 12380 9274 12436 9276
rect 12460 9274 12516 9276
rect 12220 9222 12266 9274
rect 12266 9222 12276 9274
rect 12300 9222 12330 9274
rect 12330 9222 12342 9274
rect 12342 9222 12356 9274
rect 12380 9222 12394 9274
rect 12394 9222 12406 9274
rect 12406 9222 12436 9274
rect 12460 9222 12470 9274
rect 12470 9222 12516 9274
rect 12220 9220 12276 9222
rect 12300 9220 12356 9222
rect 12380 9220 12436 9222
rect 12460 9220 12516 9222
rect 12220 8186 12276 8188
rect 12300 8186 12356 8188
rect 12380 8186 12436 8188
rect 12460 8186 12516 8188
rect 12220 8134 12266 8186
rect 12266 8134 12276 8186
rect 12300 8134 12330 8186
rect 12330 8134 12342 8186
rect 12342 8134 12356 8186
rect 12380 8134 12394 8186
rect 12394 8134 12406 8186
rect 12406 8134 12436 8186
rect 12460 8134 12470 8186
rect 12470 8134 12516 8186
rect 12220 8132 12276 8134
rect 12300 8132 12356 8134
rect 12380 8132 12436 8134
rect 12460 8132 12516 8134
rect 12220 7098 12276 7100
rect 12300 7098 12356 7100
rect 12380 7098 12436 7100
rect 12460 7098 12516 7100
rect 12220 7046 12266 7098
rect 12266 7046 12276 7098
rect 12300 7046 12330 7098
rect 12330 7046 12342 7098
rect 12342 7046 12356 7098
rect 12380 7046 12394 7098
rect 12394 7046 12406 7098
rect 12406 7046 12436 7098
rect 12460 7046 12470 7098
rect 12470 7046 12516 7098
rect 12220 7044 12276 7046
rect 12300 7044 12356 7046
rect 12380 7044 12436 7046
rect 12460 7044 12516 7046
rect 12220 6010 12276 6012
rect 12300 6010 12356 6012
rect 12380 6010 12436 6012
rect 12460 6010 12516 6012
rect 12220 5958 12266 6010
rect 12266 5958 12276 6010
rect 12300 5958 12330 6010
rect 12330 5958 12342 6010
rect 12342 5958 12356 6010
rect 12380 5958 12394 6010
rect 12394 5958 12406 6010
rect 12406 5958 12436 6010
rect 12460 5958 12470 6010
rect 12470 5958 12516 6010
rect 12220 5956 12276 5958
rect 12300 5956 12356 5958
rect 12380 5956 12436 5958
rect 12460 5956 12516 5958
rect 11426 5652 11428 5672
rect 11428 5652 11480 5672
rect 11480 5652 11482 5672
rect 11426 5616 11482 5652
rect 12220 4922 12276 4924
rect 12300 4922 12356 4924
rect 12380 4922 12436 4924
rect 12460 4922 12516 4924
rect 12220 4870 12266 4922
rect 12266 4870 12276 4922
rect 12300 4870 12330 4922
rect 12330 4870 12342 4922
rect 12342 4870 12356 4922
rect 12380 4870 12394 4922
rect 12394 4870 12406 4922
rect 12406 4870 12436 4922
rect 12460 4870 12470 4922
rect 12470 4870 12516 4922
rect 12220 4868 12276 4870
rect 12300 4868 12356 4870
rect 12380 4868 12436 4870
rect 12460 4868 12516 4870
rect 12220 3834 12276 3836
rect 12300 3834 12356 3836
rect 12380 3834 12436 3836
rect 12460 3834 12516 3836
rect 12220 3782 12266 3834
rect 12266 3782 12276 3834
rect 12300 3782 12330 3834
rect 12330 3782 12342 3834
rect 12342 3782 12356 3834
rect 12380 3782 12394 3834
rect 12394 3782 12406 3834
rect 12406 3782 12436 3834
rect 12460 3782 12470 3834
rect 12470 3782 12516 3834
rect 12220 3780 12276 3782
rect 12300 3780 12356 3782
rect 12380 3780 12436 3782
rect 12460 3780 12516 3782
rect 12220 2746 12276 2748
rect 12300 2746 12356 2748
rect 12380 2746 12436 2748
rect 12460 2746 12516 2748
rect 12220 2694 12266 2746
rect 12266 2694 12276 2746
rect 12300 2694 12330 2746
rect 12330 2694 12342 2746
rect 12342 2694 12356 2746
rect 12380 2694 12394 2746
rect 12394 2694 12406 2746
rect 12406 2694 12436 2746
rect 12460 2694 12470 2746
rect 12470 2694 12516 2746
rect 12220 2692 12276 2694
rect 12300 2692 12356 2694
rect 12380 2692 12436 2694
rect 12460 2692 12516 2694
rect 12220 1658 12276 1660
rect 12300 1658 12356 1660
rect 12380 1658 12436 1660
rect 12460 1658 12516 1660
rect 12220 1606 12266 1658
rect 12266 1606 12276 1658
rect 12300 1606 12330 1658
rect 12330 1606 12342 1658
rect 12342 1606 12356 1658
rect 12380 1606 12394 1658
rect 12394 1606 12406 1658
rect 12406 1606 12436 1658
rect 12460 1606 12470 1658
rect 12470 1606 12516 1658
rect 12220 1604 12276 1606
rect 12300 1604 12356 1606
rect 12380 1604 12436 1606
rect 12460 1604 12516 1606
rect 16220 17434 16276 17436
rect 16300 17434 16356 17436
rect 16380 17434 16436 17436
rect 16460 17434 16516 17436
rect 16220 17382 16266 17434
rect 16266 17382 16276 17434
rect 16300 17382 16330 17434
rect 16330 17382 16342 17434
rect 16342 17382 16356 17434
rect 16380 17382 16394 17434
rect 16394 17382 16406 17434
rect 16406 17382 16436 17434
rect 16460 17382 16470 17434
rect 16470 17382 16516 17434
rect 16220 17380 16276 17382
rect 16300 17380 16356 17382
rect 16380 17380 16436 17382
rect 16460 17380 16516 17382
rect 16220 16346 16276 16348
rect 16300 16346 16356 16348
rect 16380 16346 16436 16348
rect 16460 16346 16516 16348
rect 16220 16294 16266 16346
rect 16266 16294 16276 16346
rect 16300 16294 16330 16346
rect 16330 16294 16342 16346
rect 16342 16294 16356 16346
rect 16380 16294 16394 16346
rect 16394 16294 16406 16346
rect 16406 16294 16436 16346
rect 16460 16294 16470 16346
rect 16470 16294 16516 16346
rect 16220 16292 16276 16294
rect 16300 16292 16356 16294
rect 16380 16292 16436 16294
rect 16460 16292 16516 16294
rect 17038 16088 17094 16144
rect 20220 20154 20276 20156
rect 20300 20154 20356 20156
rect 20380 20154 20436 20156
rect 20460 20154 20516 20156
rect 20220 20102 20266 20154
rect 20266 20102 20276 20154
rect 20300 20102 20330 20154
rect 20330 20102 20342 20154
rect 20342 20102 20356 20154
rect 20380 20102 20394 20154
rect 20394 20102 20406 20154
rect 20406 20102 20436 20154
rect 20460 20102 20470 20154
rect 20470 20102 20516 20154
rect 20220 20100 20276 20102
rect 20300 20100 20356 20102
rect 20380 20100 20436 20102
rect 20460 20100 20516 20102
rect 20220 19066 20276 19068
rect 20300 19066 20356 19068
rect 20380 19066 20436 19068
rect 20460 19066 20516 19068
rect 20220 19014 20266 19066
rect 20266 19014 20276 19066
rect 20300 19014 20330 19066
rect 20330 19014 20342 19066
rect 20342 19014 20356 19066
rect 20380 19014 20394 19066
rect 20394 19014 20406 19066
rect 20406 19014 20436 19066
rect 20460 19014 20470 19066
rect 20470 19014 20516 19066
rect 20220 19012 20276 19014
rect 20300 19012 20356 19014
rect 20380 19012 20436 19014
rect 20460 19012 20516 19014
rect 20220 17978 20276 17980
rect 20300 17978 20356 17980
rect 20380 17978 20436 17980
rect 20460 17978 20516 17980
rect 20220 17926 20266 17978
rect 20266 17926 20276 17978
rect 20300 17926 20330 17978
rect 20330 17926 20342 17978
rect 20342 17926 20356 17978
rect 20380 17926 20394 17978
rect 20394 17926 20406 17978
rect 20406 17926 20436 17978
rect 20460 17926 20470 17978
rect 20470 17926 20516 17978
rect 20220 17924 20276 17926
rect 20300 17924 20356 17926
rect 20380 17924 20436 17926
rect 20460 17924 20516 17926
rect 20220 16890 20276 16892
rect 20300 16890 20356 16892
rect 20380 16890 20436 16892
rect 20460 16890 20516 16892
rect 20220 16838 20266 16890
rect 20266 16838 20276 16890
rect 20300 16838 20330 16890
rect 20330 16838 20342 16890
rect 20342 16838 20356 16890
rect 20380 16838 20394 16890
rect 20394 16838 20406 16890
rect 20406 16838 20436 16890
rect 20460 16838 20470 16890
rect 20470 16838 20516 16890
rect 20220 16836 20276 16838
rect 20300 16836 20356 16838
rect 20380 16836 20436 16838
rect 20460 16836 20516 16838
rect 24220 20698 24276 20700
rect 24300 20698 24356 20700
rect 24380 20698 24436 20700
rect 24460 20698 24516 20700
rect 24220 20646 24266 20698
rect 24266 20646 24276 20698
rect 24300 20646 24330 20698
rect 24330 20646 24342 20698
rect 24342 20646 24356 20698
rect 24380 20646 24394 20698
rect 24394 20646 24406 20698
rect 24406 20646 24436 20698
rect 24460 20646 24470 20698
rect 24470 20646 24516 20698
rect 24220 20644 24276 20646
rect 24300 20644 24356 20646
rect 24380 20644 24436 20646
rect 24460 20644 24516 20646
rect 24858 19624 24914 19680
rect 24220 19610 24276 19612
rect 24300 19610 24356 19612
rect 24380 19610 24436 19612
rect 24460 19610 24516 19612
rect 24220 19558 24266 19610
rect 24266 19558 24276 19610
rect 24300 19558 24330 19610
rect 24330 19558 24342 19610
rect 24342 19558 24356 19610
rect 24380 19558 24394 19610
rect 24394 19558 24406 19610
rect 24406 19558 24436 19610
rect 24460 19558 24470 19610
rect 24470 19558 24516 19610
rect 24220 19556 24276 19558
rect 24300 19556 24356 19558
rect 24380 19556 24436 19558
rect 24460 19556 24516 19558
rect 24220 18522 24276 18524
rect 24300 18522 24356 18524
rect 24380 18522 24436 18524
rect 24460 18522 24516 18524
rect 24220 18470 24266 18522
rect 24266 18470 24276 18522
rect 24300 18470 24330 18522
rect 24330 18470 24342 18522
rect 24342 18470 24356 18522
rect 24380 18470 24394 18522
rect 24394 18470 24406 18522
rect 24406 18470 24436 18522
rect 24460 18470 24470 18522
rect 24470 18470 24516 18522
rect 24220 18468 24276 18470
rect 24300 18468 24356 18470
rect 24380 18468 24436 18470
rect 24460 18468 24516 18470
rect 24220 17434 24276 17436
rect 24300 17434 24356 17436
rect 24380 17434 24436 17436
rect 24460 17434 24516 17436
rect 24220 17382 24266 17434
rect 24266 17382 24276 17434
rect 24300 17382 24330 17434
rect 24330 17382 24342 17434
rect 24342 17382 24356 17434
rect 24380 17382 24394 17434
rect 24394 17382 24406 17434
rect 24406 17382 24436 17434
rect 24460 17382 24470 17434
rect 24470 17382 24516 17434
rect 24220 17380 24276 17382
rect 24300 17380 24356 17382
rect 24380 17380 24436 17382
rect 24460 17380 24516 17382
rect 24220 16346 24276 16348
rect 24300 16346 24356 16348
rect 24380 16346 24436 16348
rect 24460 16346 24516 16348
rect 24220 16294 24266 16346
rect 24266 16294 24276 16346
rect 24300 16294 24330 16346
rect 24330 16294 24342 16346
rect 24342 16294 24356 16346
rect 24380 16294 24394 16346
rect 24394 16294 24406 16346
rect 24406 16294 24436 16346
rect 24460 16294 24470 16346
rect 24470 16294 24516 16346
rect 24220 16292 24276 16294
rect 24300 16292 24356 16294
rect 24380 16292 24436 16294
rect 24460 16292 24516 16294
rect 24858 16088 24914 16144
rect 20220 15802 20276 15804
rect 20300 15802 20356 15804
rect 20380 15802 20436 15804
rect 20460 15802 20516 15804
rect 20220 15750 20266 15802
rect 20266 15750 20276 15802
rect 20300 15750 20330 15802
rect 20330 15750 20342 15802
rect 20342 15750 20356 15802
rect 20380 15750 20394 15802
rect 20394 15750 20406 15802
rect 20406 15750 20436 15802
rect 20460 15750 20470 15802
rect 20470 15750 20516 15802
rect 20220 15748 20276 15750
rect 20300 15748 20356 15750
rect 20380 15748 20436 15750
rect 20460 15748 20516 15750
rect 16220 15258 16276 15260
rect 16300 15258 16356 15260
rect 16380 15258 16436 15260
rect 16460 15258 16516 15260
rect 16220 15206 16266 15258
rect 16266 15206 16276 15258
rect 16300 15206 16330 15258
rect 16330 15206 16342 15258
rect 16342 15206 16356 15258
rect 16380 15206 16394 15258
rect 16394 15206 16406 15258
rect 16406 15206 16436 15258
rect 16460 15206 16470 15258
rect 16470 15206 16516 15258
rect 16220 15204 16276 15206
rect 16300 15204 16356 15206
rect 16380 15204 16436 15206
rect 16460 15204 16516 15206
rect 24220 15258 24276 15260
rect 24300 15258 24356 15260
rect 24380 15258 24436 15260
rect 24460 15258 24516 15260
rect 24220 15206 24266 15258
rect 24266 15206 24276 15258
rect 24300 15206 24330 15258
rect 24330 15206 24342 15258
rect 24342 15206 24356 15258
rect 24380 15206 24394 15258
rect 24394 15206 24406 15258
rect 24406 15206 24436 15258
rect 24460 15206 24470 15258
rect 24470 15206 24516 15258
rect 24220 15204 24276 15206
rect 24300 15204 24356 15206
rect 24380 15204 24436 15206
rect 24460 15204 24516 15206
rect 16220 14170 16276 14172
rect 16300 14170 16356 14172
rect 16380 14170 16436 14172
rect 16460 14170 16516 14172
rect 16220 14118 16266 14170
rect 16266 14118 16276 14170
rect 16300 14118 16330 14170
rect 16330 14118 16342 14170
rect 16342 14118 16356 14170
rect 16380 14118 16394 14170
rect 16394 14118 16406 14170
rect 16406 14118 16436 14170
rect 16460 14118 16470 14170
rect 16470 14118 16516 14170
rect 16220 14116 16276 14118
rect 16300 14116 16356 14118
rect 16380 14116 16436 14118
rect 16460 14116 16516 14118
rect 20220 14714 20276 14716
rect 20300 14714 20356 14716
rect 20380 14714 20436 14716
rect 20460 14714 20516 14716
rect 20220 14662 20266 14714
rect 20266 14662 20276 14714
rect 20300 14662 20330 14714
rect 20330 14662 20342 14714
rect 20342 14662 20356 14714
rect 20380 14662 20394 14714
rect 20394 14662 20406 14714
rect 20406 14662 20436 14714
rect 20460 14662 20470 14714
rect 20470 14662 20516 14714
rect 20220 14660 20276 14662
rect 20300 14660 20356 14662
rect 20380 14660 20436 14662
rect 20460 14660 20516 14662
rect 24220 14170 24276 14172
rect 24300 14170 24356 14172
rect 24380 14170 24436 14172
rect 24460 14170 24516 14172
rect 24220 14118 24266 14170
rect 24266 14118 24276 14170
rect 24300 14118 24330 14170
rect 24330 14118 24342 14170
rect 24342 14118 24356 14170
rect 24380 14118 24394 14170
rect 24394 14118 24406 14170
rect 24406 14118 24436 14170
rect 24460 14118 24470 14170
rect 24470 14118 24516 14170
rect 24220 14116 24276 14118
rect 24300 14116 24356 14118
rect 24380 14116 24436 14118
rect 24460 14116 24516 14118
rect 16220 13082 16276 13084
rect 16300 13082 16356 13084
rect 16380 13082 16436 13084
rect 16460 13082 16516 13084
rect 16220 13030 16266 13082
rect 16266 13030 16276 13082
rect 16300 13030 16330 13082
rect 16330 13030 16342 13082
rect 16342 13030 16356 13082
rect 16380 13030 16394 13082
rect 16394 13030 16406 13082
rect 16406 13030 16436 13082
rect 16460 13030 16470 13082
rect 16470 13030 16516 13082
rect 16220 13028 16276 13030
rect 16300 13028 16356 13030
rect 16380 13028 16436 13030
rect 16460 13028 16516 13030
rect 16220 11994 16276 11996
rect 16300 11994 16356 11996
rect 16380 11994 16436 11996
rect 16460 11994 16516 11996
rect 16220 11942 16266 11994
rect 16266 11942 16276 11994
rect 16300 11942 16330 11994
rect 16330 11942 16342 11994
rect 16342 11942 16356 11994
rect 16380 11942 16394 11994
rect 16394 11942 16406 11994
rect 16406 11942 16436 11994
rect 16460 11942 16470 11994
rect 16470 11942 16516 11994
rect 16220 11940 16276 11942
rect 16300 11940 16356 11942
rect 16380 11940 16436 11942
rect 16460 11940 16516 11942
rect 16220 10906 16276 10908
rect 16300 10906 16356 10908
rect 16380 10906 16436 10908
rect 16460 10906 16516 10908
rect 16220 10854 16266 10906
rect 16266 10854 16276 10906
rect 16300 10854 16330 10906
rect 16330 10854 16342 10906
rect 16342 10854 16356 10906
rect 16380 10854 16394 10906
rect 16394 10854 16406 10906
rect 16406 10854 16436 10906
rect 16460 10854 16470 10906
rect 16470 10854 16516 10906
rect 16220 10852 16276 10854
rect 16300 10852 16356 10854
rect 16380 10852 16436 10854
rect 16460 10852 16516 10854
rect 20220 13626 20276 13628
rect 20300 13626 20356 13628
rect 20380 13626 20436 13628
rect 20460 13626 20516 13628
rect 20220 13574 20266 13626
rect 20266 13574 20276 13626
rect 20300 13574 20330 13626
rect 20330 13574 20342 13626
rect 20342 13574 20356 13626
rect 20380 13574 20394 13626
rect 20394 13574 20406 13626
rect 20406 13574 20436 13626
rect 20460 13574 20470 13626
rect 20470 13574 20516 13626
rect 20220 13572 20276 13574
rect 20300 13572 20356 13574
rect 20380 13572 20436 13574
rect 20460 13572 20516 13574
rect 24220 13082 24276 13084
rect 24300 13082 24356 13084
rect 24380 13082 24436 13084
rect 24460 13082 24516 13084
rect 24220 13030 24266 13082
rect 24266 13030 24276 13082
rect 24300 13030 24330 13082
rect 24330 13030 24342 13082
rect 24342 13030 24356 13082
rect 24380 13030 24394 13082
rect 24394 13030 24406 13082
rect 24406 13030 24436 13082
rect 24460 13030 24470 13082
rect 24470 13030 24516 13082
rect 24220 13028 24276 13030
rect 24300 13028 24356 13030
rect 24380 13028 24436 13030
rect 24460 13028 24516 13030
rect 24950 12552 25006 12608
rect 20220 12538 20276 12540
rect 20300 12538 20356 12540
rect 20380 12538 20436 12540
rect 20460 12538 20516 12540
rect 20220 12486 20266 12538
rect 20266 12486 20276 12538
rect 20300 12486 20330 12538
rect 20330 12486 20342 12538
rect 20342 12486 20356 12538
rect 20380 12486 20394 12538
rect 20394 12486 20406 12538
rect 20406 12486 20436 12538
rect 20460 12486 20470 12538
rect 20470 12486 20516 12538
rect 20220 12484 20276 12486
rect 20300 12484 20356 12486
rect 20380 12484 20436 12486
rect 20460 12484 20516 12486
rect 16220 9818 16276 9820
rect 16300 9818 16356 9820
rect 16380 9818 16436 9820
rect 16460 9818 16516 9820
rect 16220 9766 16266 9818
rect 16266 9766 16276 9818
rect 16300 9766 16330 9818
rect 16330 9766 16342 9818
rect 16342 9766 16356 9818
rect 16380 9766 16394 9818
rect 16394 9766 16406 9818
rect 16406 9766 16436 9818
rect 16460 9766 16470 9818
rect 16470 9766 16516 9818
rect 16220 9764 16276 9766
rect 16300 9764 16356 9766
rect 16380 9764 16436 9766
rect 16460 9764 16516 9766
rect 15934 9016 15990 9072
rect 16220 8730 16276 8732
rect 16300 8730 16356 8732
rect 16380 8730 16436 8732
rect 16460 8730 16516 8732
rect 16220 8678 16266 8730
rect 16266 8678 16276 8730
rect 16300 8678 16330 8730
rect 16330 8678 16342 8730
rect 16342 8678 16356 8730
rect 16380 8678 16394 8730
rect 16394 8678 16406 8730
rect 16406 8678 16436 8730
rect 16460 8678 16470 8730
rect 16470 8678 16516 8730
rect 16220 8676 16276 8678
rect 16300 8676 16356 8678
rect 16380 8676 16436 8678
rect 16460 8676 16516 8678
rect 16220 7642 16276 7644
rect 16300 7642 16356 7644
rect 16380 7642 16436 7644
rect 16460 7642 16516 7644
rect 16220 7590 16266 7642
rect 16266 7590 16276 7642
rect 16300 7590 16330 7642
rect 16330 7590 16342 7642
rect 16342 7590 16356 7642
rect 16380 7590 16394 7642
rect 16394 7590 16406 7642
rect 16406 7590 16436 7642
rect 16460 7590 16470 7642
rect 16470 7590 16516 7642
rect 16220 7588 16276 7590
rect 16300 7588 16356 7590
rect 16380 7588 16436 7590
rect 16460 7588 16516 7590
rect 16220 6554 16276 6556
rect 16300 6554 16356 6556
rect 16380 6554 16436 6556
rect 16460 6554 16516 6556
rect 16220 6502 16266 6554
rect 16266 6502 16276 6554
rect 16300 6502 16330 6554
rect 16330 6502 16342 6554
rect 16342 6502 16356 6554
rect 16380 6502 16394 6554
rect 16394 6502 16406 6554
rect 16406 6502 16436 6554
rect 16460 6502 16470 6554
rect 16470 6502 16516 6554
rect 16220 6500 16276 6502
rect 16300 6500 16356 6502
rect 16380 6500 16436 6502
rect 16460 6500 16516 6502
rect 15750 5616 15806 5672
rect 16220 5466 16276 5468
rect 16300 5466 16356 5468
rect 16380 5466 16436 5468
rect 16460 5466 16516 5468
rect 16220 5414 16266 5466
rect 16266 5414 16276 5466
rect 16300 5414 16330 5466
rect 16330 5414 16342 5466
rect 16342 5414 16356 5466
rect 16380 5414 16394 5466
rect 16394 5414 16406 5466
rect 16406 5414 16436 5466
rect 16460 5414 16470 5466
rect 16470 5414 16516 5466
rect 16220 5412 16276 5414
rect 16300 5412 16356 5414
rect 16380 5412 16436 5414
rect 16460 5412 16516 5414
rect 16220 4378 16276 4380
rect 16300 4378 16356 4380
rect 16380 4378 16436 4380
rect 16460 4378 16516 4380
rect 16220 4326 16266 4378
rect 16266 4326 16276 4378
rect 16300 4326 16330 4378
rect 16330 4326 16342 4378
rect 16342 4326 16356 4378
rect 16380 4326 16394 4378
rect 16394 4326 16406 4378
rect 16406 4326 16436 4378
rect 16460 4326 16470 4378
rect 16470 4326 16516 4378
rect 16220 4324 16276 4326
rect 16300 4324 16356 4326
rect 16380 4324 16436 4326
rect 16460 4324 16516 4326
rect 16220 3290 16276 3292
rect 16300 3290 16356 3292
rect 16380 3290 16436 3292
rect 16460 3290 16516 3292
rect 16220 3238 16266 3290
rect 16266 3238 16276 3290
rect 16300 3238 16330 3290
rect 16330 3238 16342 3290
rect 16342 3238 16356 3290
rect 16380 3238 16394 3290
rect 16394 3238 16406 3290
rect 16406 3238 16436 3290
rect 16460 3238 16470 3290
rect 16470 3238 16516 3290
rect 16220 3236 16276 3238
rect 16300 3236 16356 3238
rect 16380 3236 16436 3238
rect 16460 3236 16516 3238
rect 24220 11994 24276 11996
rect 24300 11994 24356 11996
rect 24380 11994 24436 11996
rect 24460 11994 24516 11996
rect 24220 11942 24266 11994
rect 24266 11942 24276 11994
rect 24300 11942 24330 11994
rect 24330 11942 24342 11994
rect 24342 11942 24356 11994
rect 24380 11942 24394 11994
rect 24394 11942 24406 11994
rect 24406 11942 24436 11994
rect 24460 11942 24470 11994
rect 24470 11942 24516 11994
rect 24220 11940 24276 11942
rect 24300 11940 24356 11942
rect 24380 11940 24436 11942
rect 24460 11940 24516 11942
rect 20220 11450 20276 11452
rect 20300 11450 20356 11452
rect 20380 11450 20436 11452
rect 20460 11450 20516 11452
rect 20220 11398 20266 11450
rect 20266 11398 20276 11450
rect 20300 11398 20330 11450
rect 20330 11398 20342 11450
rect 20342 11398 20356 11450
rect 20380 11398 20394 11450
rect 20394 11398 20406 11450
rect 20406 11398 20436 11450
rect 20460 11398 20470 11450
rect 20470 11398 20516 11450
rect 20220 11396 20276 11398
rect 20300 11396 20356 11398
rect 20380 11396 20436 11398
rect 20460 11396 20516 11398
rect 20220 10362 20276 10364
rect 20300 10362 20356 10364
rect 20380 10362 20436 10364
rect 20460 10362 20516 10364
rect 20220 10310 20266 10362
rect 20266 10310 20276 10362
rect 20300 10310 20330 10362
rect 20330 10310 20342 10362
rect 20342 10310 20356 10362
rect 20380 10310 20394 10362
rect 20394 10310 20406 10362
rect 20406 10310 20436 10362
rect 20460 10310 20470 10362
rect 20470 10310 20516 10362
rect 20220 10308 20276 10310
rect 20300 10308 20356 10310
rect 20380 10308 20436 10310
rect 20460 10308 20516 10310
rect 20220 9274 20276 9276
rect 20300 9274 20356 9276
rect 20380 9274 20436 9276
rect 20460 9274 20516 9276
rect 20220 9222 20266 9274
rect 20266 9222 20276 9274
rect 20300 9222 20330 9274
rect 20330 9222 20342 9274
rect 20342 9222 20356 9274
rect 20380 9222 20394 9274
rect 20394 9222 20406 9274
rect 20406 9222 20436 9274
rect 20460 9222 20470 9274
rect 20470 9222 20516 9274
rect 20220 9220 20276 9222
rect 20300 9220 20356 9222
rect 20380 9220 20436 9222
rect 20460 9220 20516 9222
rect 24220 10906 24276 10908
rect 24300 10906 24356 10908
rect 24380 10906 24436 10908
rect 24460 10906 24516 10908
rect 24220 10854 24266 10906
rect 24266 10854 24276 10906
rect 24300 10854 24330 10906
rect 24330 10854 24342 10906
rect 24342 10854 24356 10906
rect 24380 10854 24394 10906
rect 24394 10854 24406 10906
rect 24406 10854 24436 10906
rect 24460 10854 24470 10906
rect 24470 10854 24516 10906
rect 24220 10852 24276 10854
rect 24300 10852 24356 10854
rect 24380 10852 24436 10854
rect 24460 10852 24516 10854
rect 20220 8186 20276 8188
rect 20300 8186 20356 8188
rect 20380 8186 20436 8188
rect 20460 8186 20516 8188
rect 20220 8134 20266 8186
rect 20266 8134 20276 8186
rect 20300 8134 20330 8186
rect 20330 8134 20342 8186
rect 20342 8134 20356 8186
rect 20380 8134 20394 8186
rect 20394 8134 20406 8186
rect 20406 8134 20436 8186
rect 20460 8134 20470 8186
rect 20470 8134 20516 8186
rect 20220 8132 20276 8134
rect 20300 8132 20356 8134
rect 20380 8132 20436 8134
rect 20460 8132 20516 8134
rect 20220 7098 20276 7100
rect 20300 7098 20356 7100
rect 20380 7098 20436 7100
rect 20460 7098 20516 7100
rect 20220 7046 20266 7098
rect 20266 7046 20276 7098
rect 20300 7046 20330 7098
rect 20330 7046 20342 7098
rect 20342 7046 20356 7098
rect 20380 7046 20394 7098
rect 20394 7046 20406 7098
rect 20406 7046 20436 7098
rect 20460 7046 20470 7098
rect 20470 7046 20516 7098
rect 20220 7044 20276 7046
rect 20300 7044 20356 7046
rect 20380 7044 20436 7046
rect 20460 7044 20516 7046
rect 20220 6010 20276 6012
rect 20300 6010 20356 6012
rect 20380 6010 20436 6012
rect 20460 6010 20516 6012
rect 20220 5958 20266 6010
rect 20266 5958 20276 6010
rect 20300 5958 20330 6010
rect 20330 5958 20342 6010
rect 20342 5958 20356 6010
rect 20380 5958 20394 6010
rect 20394 5958 20406 6010
rect 20406 5958 20436 6010
rect 20460 5958 20470 6010
rect 20470 5958 20516 6010
rect 20220 5956 20276 5958
rect 20300 5956 20356 5958
rect 20380 5956 20436 5958
rect 20460 5956 20516 5958
rect 16220 2202 16276 2204
rect 16300 2202 16356 2204
rect 16380 2202 16436 2204
rect 16460 2202 16516 2204
rect 16220 2150 16266 2202
rect 16266 2150 16276 2202
rect 16300 2150 16330 2202
rect 16330 2150 16342 2202
rect 16342 2150 16356 2202
rect 16380 2150 16394 2202
rect 16394 2150 16406 2202
rect 16406 2150 16436 2202
rect 16460 2150 16470 2202
rect 16470 2150 16516 2202
rect 16220 2148 16276 2150
rect 16300 2148 16356 2150
rect 16380 2148 16436 2150
rect 16460 2148 16516 2150
rect 20220 4922 20276 4924
rect 20300 4922 20356 4924
rect 20380 4922 20436 4924
rect 20460 4922 20516 4924
rect 20220 4870 20266 4922
rect 20266 4870 20276 4922
rect 20300 4870 20330 4922
rect 20330 4870 20342 4922
rect 20342 4870 20356 4922
rect 20380 4870 20394 4922
rect 20394 4870 20406 4922
rect 20406 4870 20436 4922
rect 20460 4870 20470 4922
rect 20470 4870 20516 4922
rect 20220 4868 20276 4870
rect 20300 4868 20356 4870
rect 20380 4868 20436 4870
rect 20460 4868 20516 4870
rect 20220 3834 20276 3836
rect 20300 3834 20356 3836
rect 20380 3834 20436 3836
rect 20460 3834 20516 3836
rect 20220 3782 20266 3834
rect 20266 3782 20276 3834
rect 20300 3782 20330 3834
rect 20330 3782 20342 3834
rect 20342 3782 20356 3834
rect 20380 3782 20394 3834
rect 20394 3782 20406 3834
rect 20406 3782 20436 3834
rect 20460 3782 20470 3834
rect 20470 3782 20516 3834
rect 20220 3780 20276 3782
rect 20300 3780 20356 3782
rect 20380 3780 20436 3782
rect 20460 3780 20516 3782
rect 20220 2746 20276 2748
rect 20300 2746 20356 2748
rect 20380 2746 20436 2748
rect 20460 2746 20516 2748
rect 20220 2694 20266 2746
rect 20266 2694 20276 2746
rect 20300 2694 20330 2746
rect 20330 2694 20342 2746
rect 20342 2694 20356 2746
rect 20380 2694 20394 2746
rect 20394 2694 20406 2746
rect 20406 2694 20436 2746
rect 20460 2694 20470 2746
rect 20470 2694 20516 2746
rect 20220 2692 20276 2694
rect 20300 2692 20356 2694
rect 20380 2692 20436 2694
rect 20460 2692 20516 2694
rect 24220 9818 24276 9820
rect 24300 9818 24356 9820
rect 24380 9818 24436 9820
rect 24460 9818 24516 9820
rect 24220 9766 24266 9818
rect 24266 9766 24276 9818
rect 24300 9766 24330 9818
rect 24330 9766 24342 9818
rect 24342 9766 24356 9818
rect 24380 9766 24394 9818
rect 24394 9766 24406 9818
rect 24406 9766 24436 9818
rect 24460 9766 24470 9818
rect 24470 9766 24516 9818
rect 24220 9764 24276 9766
rect 24300 9764 24356 9766
rect 24380 9764 24436 9766
rect 24460 9764 24516 9766
rect 24220 8730 24276 8732
rect 24300 8730 24356 8732
rect 24380 8730 24436 8732
rect 24460 8730 24516 8732
rect 24220 8678 24266 8730
rect 24266 8678 24276 8730
rect 24300 8678 24330 8730
rect 24330 8678 24342 8730
rect 24342 8678 24356 8730
rect 24380 8678 24394 8730
rect 24394 8678 24406 8730
rect 24406 8678 24436 8730
rect 24460 8678 24470 8730
rect 24470 8678 24516 8730
rect 24220 8676 24276 8678
rect 24300 8676 24356 8678
rect 24380 8676 24436 8678
rect 24460 8676 24516 8678
rect 24220 7642 24276 7644
rect 24300 7642 24356 7644
rect 24380 7642 24436 7644
rect 24460 7642 24516 7644
rect 24220 7590 24266 7642
rect 24266 7590 24276 7642
rect 24300 7590 24330 7642
rect 24330 7590 24342 7642
rect 24342 7590 24356 7642
rect 24380 7590 24394 7642
rect 24394 7590 24406 7642
rect 24406 7590 24436 7642
rect 24460 7590 24470 7642
rect 24470 7590 24516 7642
rect 24220 7588 24276 7590
rect 24300 7588 24356 7590
rect 24380 7588 24436 7590
rect 24460 7588 24516 7590
rect 24220 6554 24276 6556
rect 24300 6554 24356 6556
rect 24380 6554 24436 6556
rect 24460 6554 24516 6556
rect 24220 6502 24266 6554
rect 24266 6502 24276 6554
rect 24300 6502 24330 6554
rect 24330 6502 24342 6554
rect 24342 6502 24356 6554
rect 24380 6502 24394 6554
rect 24394 6502 24406 6554
rect 24406 6502 24436 6554
rect 24460 6502 24470 6554
rect 24470 6502 24516 6554
rect 24220 6500 24276 6502
rect 24300 6500 24356 6502
rect 24380 6500 24436 6502
rect 24460 6500 24516 6502
rect 24220 5466 24276 5468
rect 24300 5466 24356 5468
rect 24380 5466 24436 5468
rect 24460 5466 24516 5468
rect 24220 5414 24266 5466
rect 24266 5414 24276 5466
rect 24300 5414 24330 5466
rect 24330 5414 24342 5466
rect 24342 5414 24356 5466
rect 24380 5414 24394 5466
rect 24394 5414 24406 5466
rect 24406 5414 24436 5466
rect 24460 5414 24470 5466
rect 24470 5414 24516 5466
rect 24220 5412 24276 5414
rect 24300 5412 24356 5414
rect 24380 5412 24436 5414
rect 24460 5412 24516 5414
rect 26146 5480 26202 5536
rect 24220 4378 24276 4380
rect 24300 4378 24356 4380
rect 24380 4378 24436 4380
rect 24460 4378 24516 4380
rect 24220 4326 24266 4378
rect 24266 4326 24276 4378
rect 24300 4326 24330 4378
rect 24330 4326 24342 4378
rect 24342 4326 24356 4378
rect 24380 4326 24394 4378
rect 24394 4326 24406 4378
rect 24406 4326 24436 4378
rect 24460 4326 24470 4378
rect 24470 4326 24516 4378
rect 24220 4324 24276 4326
rect 24300 4324 24356 4326
rect 24380 4324 24436 4326
rect 24460 4324 24516 4326
rect 24220 3290 24276 3292
rect 24300 3290 24356 3292
rect 24380 3290 24436 3292
rect 24460 3290 24516 3292
rect 24220 3238 24266 3290
rect 24266 3238 24276 3290
rect 24300 3238 24330 3290
rect 24330 3238 24342 3290
rect 24342 3238 24356 3290
rect 24380 3238 24394 3290
rect 24394 3238 24406 3290
rect 24406 3238 24436 3290
rect 24460 3238 24470 3290
rect 24470 3238 24516 3290
rect 24220 3236 24276 3238
rect 24300 3236 24356 3238
rect 24380 3236 24436 3238
rect 24460 3236 24516 3238
rect 24220 2202 24276 2204
rect 24300 2202 24356 2204
rect 24380 2202 24436 2204
rect 24460 2202 24516 2204
rect 24220 2150 24266 2202
rect 24266 2150 24276 2202
rect 24300 2150 24330 2202
rect 24330 2150 24342 2202
rect 24342 2150 24356 2202
rect 24380 2150 24394 2202
rect 24394 2150 24406 2202
rect 24406 2150 24436 2202
rect 24460 2150 24470 2202
rect 24470 2150 24516 2202
rect 24220 2148 24276 2150
rect 24300 2148 24356 2150
rect 24380 2148 24436 2150
rect 24460 2148 24516 2150
rect 26146 1944 26202 2000
rect 20220 1658 20276 1660
rect 20300 1658 20356 1660
rect 20380 1658 20436 1660
rect 20460 1658 20516 1660
rect 20220 1606 20266 1658
rect 20266 1606 20276 1658
rect 20300 1606 20330 1658
rect 20330 1606 20342 1658
rect 20342 1606 20356 1658
rect 20380 1606 20394 1658
rect 20394 1606 20406 1658
rect 20406 1606 20436 1658
rect 20460 1606 20470 1658
rect 20470 1606 20516 1658
rect 20220 1604 20276 1606
rect 20300 1604 20356 1606
rect 20380 1604 20436 1606
rect 20460 1604 20516 1606
rect 8220 1114 8276 1116
rect 8300 1114 8356 1116
rect 8380 1114 8436 1116
rect 8460 1114 8516 1116
rect 8220 1062 8266 1114
rect 8266 1062 8276 1114
rect 8300 1062 8330 1114
rect 8330 1062 8342 1114
rect 8342 1062 8356 1114
rect 8380 1062 8394 1114
rect 8394 1062 8406 1114
rect 8406 1062 8436 1114
rect 8460 1062 8470 1114
rect 8470 1062 8516 1114
rect 8220 1060 8276 1062
rect 8300 1060 8356 1062
rect 8380 1060 8436 1062
rect 8460 1060 8516 1062
rect 16220 1114 16276 1116
rect 16300 1114 16356 1116
rect 16380 1114 16436 1116
rect 16460 1114 16516 1116
rect 16220 1062 16266 1114
rect 16266 1062 16276 1114
rect 16300 1062 16330 1114
rect 16330 1062 16342 1114
rect 16342 1062 16356 1114
rect 16380 1062 16394 1114
rect 16394 1062 16406 1114
rect 16406 1062 16436 1114
rect 16460 1062 16470 1114
rect 16470 1062 16516 1114
rect 16220 1060 16276 1062
rect 16300 1060 16356 1062
rect 16380 1060 16436 1062
rect 16460 1060 16516 1062
rect 24220 1114 24276 1116
rect 24300 1114 24356 1116
rect 24380 1114 24436 1116
rect 24460 1114 24516 1116
rect 24220 1062 24266 1114
rect 24266 1062 24276 1114
rect 24300 1062 24330 1114
rect 24330 1062 24342 1114
rect 24342 1062 24356 1114
rect 24380 1062 24394 1114
rect 24394 1062 24406 1114
rect 24406 1062 24436 1114
rect 24460 1062 24470 1114
rect 24470 1062 24516 1114
rect 24220 1060 24276 1062
rect 24300 1060 24356 1062
rect 24380 1060 24436 1062
rect 24460 1060 24516 1062
<< metal3 >>
rect 0 20770 800 20800
rect 6729 20770 6795 20773
rect 0 20768 6795 20770
rect 0 20712 6734 20768
rect 6790 20712 6795 20768
rect 0 20710 6795 20712
rect 0 20680 800 20710
rect 6729 20707 6795 20710
rect 8210 20704 8526 20705
rect 8210 20640 8216 20704
rect 8280 20640 8296 20704
rect 8360 20640 8376 20704
rect 8440 20640 8456 20704
rect 8520 20640 8526 20704
rect 8210 20639 8526 20640
rect 16210 20704 16526 20705
rect 16210 20640 16216 20704
rect 16280 20640 16296 20704
rect 16360 20640 16376 20704
rect 16440 20640 16456 20704
rect 16520 20640 16526 20704
rect 16210 20639 16526 20640
rect 24210 20704 24526 20705
rect 24210 20640 24216 20704
rect 24280 20640 24296 20704
rect 24360 20640 24376 20704
rect 24440 20640 24456 20704
rect 24520 20640 24526 20704
rect 24210 20639 24526 20640
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 12210 20160 12526 20161
rect 12210 20096 12216 20160
rect 12280 20096 12296 20160
rect 12360 20096 12376 20160
rect 12440 20096 12456 20160
rect 12520 20096 12526 20160
rect 12210 20095 12526 20096
rect 20210 20160 20526 20161
rect 20210 20096 20216 20160
rect 20280 20096 20296 20160
rect 20360 20096 20376 20160
rect 20440 20096 20456 20160
rect 20520 20096 20526 20160
rect 20210 20095 20526 20096
rect 10777 19818 10843 19821
rect 16665 19818 16731 19821
rect 10777 19816 16731 19818
rect 10777 19760 10782 19816
rect 10838 19760 16670 19816
rect 16726 19760 16731 19816
rect 10777 19758 16731 19760
rect 10777 19755 10843 19758
rect 16665 19755 16731 19758
rect 0 19682 800 19712
rect 4613 19682 4679 19685
rect 0 19680 4679 19682
rect 0 19624 4618 19680
rect 4674 19624 4679 19680
rect 0 19622 4679 19624
rect 0 19592 800 19622
rect 4613 19619 4679 19622
rect 24853 19682 24919 19685
rect 26200 19682 27000 19712
rect 24853 19680 27000 19682
rect 24853 19624 24858 19680
rect 24914 19624 27000 19680
rect 24853 19622 27000 19624
rect 24853 19619 24919 19622
rect 8210 19616 8526 19617
rect 8210 19552 8216 19616
rect 8280 19552 8296 19616
rect 8360 19552 8376 19616
rect 8440 19552 8456 19616
rect 8520 19552 8526 19616
rect 8210 19551 8526 19552
rect 16210 19616 16526 19617
rect 16210 19552 16216 19616
rect 16280 19552 16296 19616
rect 16360 19552 16376 19616
rect 16440 19552 16456 19616
rect 16520 19552 16526 19616
rect 16210 19551 16526 19552
rect 24210 19616 24526 19617
rect 24210 19552 24216 19616
rect 24280 19552 24296 19616
rect 24360 19552 24376 19616
rect 24440 19552 24456 19616
rect 24520 19552 24526 19616
rect 26200 19592 27000 19622
rect 24210 19551 24526 19552
rect 11462 19076 11468 19140
rect 11532 19138 11538 19140
rect 11605 19138 11671 19141
rect 11532 19136 11671 19138
rect 11532 19080 11610 19136
rect 11666 19080 11671 19136
rect 11532 19078 11671 19080
rect 11532 19076 11538 19078
rect 11605 19075 11671 19078
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 12210 19072 12526 19073
rect 12210 19008 12216 19072
rect 12280 19008 12296 19072
rect 12360 19008 12376 19072
rect 12440 19008 12456 19072
rect 12520 19008 12526 19072
rect 12210 19007 12526 19008
rect 20210 19072 20526 19073
rect 20210 19008 20216 19072
rect 20280 19008 20296 19072
rect 20360 19008 20376 19072
rect 20440 19008 20456 19072
rect 20520 19008 20526 19072
rect 20210 19007 20526 19008
rect 11697 18868 11763 18869
rect 11646 18866 11652 18868
rect 11606 18806 11652 18866
rect 11716 18864 11763 18868
rect 11758 18808 11763 18864
rect 11646 18804 11652 18806
rect 11716 18804 11763 18808
rect 11697 18803 11763 18804
rect 12065 18866 12131 18869
rect 12433 18866 12499 18869
rect 13813 18866 13879 18869
rect 12065 18864 13879 18866
rect 12065 18808 12070 18864
rect 12126 18808 12438 18864
rect 12494 18808 13818 18864
rect 13874 18808 13879 18864
rect 12065 18806 13879 18808
rect 12065 18803 12131 18806
rect 12433 18803 12499 18806
rect 13813 18803 13879 18806
rect 11329 18730 11395 18733
rect 12617 18730 12683 18733
rect 11329 18728 12683 18730
rect 11329 18672 11334 18728
rect 11390 18672 12622 18728
rect 12678 18672 12683 18728
rect 11329 18670 12683 18672
rect 11329 18667 11395 18670
rect 12617 18667 12683 18670
rect 0 18594 800 18624
rect 3969 18594 4035 18597
rect 0 18592 4035 18594
rect 0 18536 3974 18592
rect 4030 18536 4035 18592
rect 0 18534 4035 18536
rect 0 18504 800 18534
rect 3969 18531 4035 18534
rect 11421 18594 11487 18597
rect 15469 18594 15535 18597
rect 11421 18592 15535 18594
rect 11421 18536 11426 18592
rect 11482 18536 15474 18592
rect 15530 18536 15535 18592
rect 11421 18534 15535 18536
rect 11421 18531 11487 18534
rect 15469 18531 15535 18534
rect 8210 18528 8526 18529
rect 8210 18464 8216 18528
rect 8280 18464 8296 18528
rect 8360 18464 8376 18528
rect 8440 18464 8456 18528
rect 8520 18464 8526 18528
rect 8210 18463 8526 18464
rect 16210 18528 16526 18529
rect 16210 18464 16216 18528
rect 16280 18464 16296 18528
rect 16360 18464 16376 18528
rect 16440 18464 16456 18528
rect 16520 18464 16526 18528
rect 16210 18463 16526 18464
rect 24210 18528 24526 18529
rect 24210 18464 24216 18528
rect 24280 18464 24296 18528
rect 24360 18464 24376 18528
rect 24440 18464 24456 18528
rect 24520 18464 24526 18528
rect 24210 18463 24526 18464
rect 11421 18458 11487 18461
rect 12341 18458 12407 18461
rect 11421 18456 12407 18458
rect 11421 18400 11426 18456
rect 11482 18400 12346 18456
rect 12402 18400 12407 18456
rect 11421 18398 12407 18400
rect 11421 18395 11487 18398
rect 12341 18395 12407 18398
rect 10961 18322 11027 18325
rect 12709 18322 12775 18325
rect 13445 18322 13511 18325
rect 10961 18320 13511 18322
rect 10961 18264 10966 18320
rect 11022 18264 12714 18320
rect 12770 18264 13450 18320
rect 13506 18264 13511 18320
rect 10961 18262 13511 18264
rect 10961 18259 11027 18262
rect 12709 18259 12775 18262
rect 13445 18259 13511 18262
rect 10409 18186 10475 18189
rect 12065 18186 12131 18189
rect 10409 18184 12131 18186
rect 10409 18128 10414 18184
rect 10470 18128 12070 18184
rect 12126 18128 12131 18184
rect 10409 18126 12131 18128
rect 10409 18123 10475 18126
rect 12065 18123 12131 18126
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 12210 17984 12526 17985
rect 12210 17920 12216 17984
rect 12280 17920 12296 17984
rect 12360 17920 12376 17984
rect 12440 17920 12456 17984
rect 12520 17920 12526 17984
rect 12210 17919 12526 17920
rect 20210 17984 20526 17985
rect 20210 17920 20216 17984
rect 20280 17920 20296 17984
rect 20360 17920 20376 17984
rect 20440 17920 20456 17984
rect 20520 17920 20526 17984
rect 20210 17919 20526 17920
rect 11462 17852 11468 17916
rect 11532 17914 11538 17916
rect 11605 17914 11671 17917
rect 11532 17912 11671 17914
rect 11532 17856 11610 17912
rect 11666 17856 11671 17912
rect 11532 17854 11671 17856
rect 11532 17852 11538 17854
rect 11605 17851 11671 17854
rect 10869 17778 10935 17781
rect 12893 17778 12959 17781
rect 10869 17776 12959 17778
rect 10869 17720 10874 17776
rect 10930 17720 12898 17776
rect 12954 17720 12959 17776
rect 10869 17718 12959 17720
rect 10869 17715 10935 17718
rect 12893 17715 12959 17718
rect 10685 17642 10751 17645
rect 13813 17642 13879 17645
rect 10685 17640 13879 17642
rect 10685 17584 10690 17640
rect 10746 17584 13818 17640
rect 13874 17584 13879 17640
rect 10685 17582 13879 17584
rect 10685 17579 10751 17582
rect 13813 17579 13879 17582
rect 0 17506 800 17536
rect 5625 17506 5691 17509
rect 0 17504 5691 17506
rect 0 17448 5630 17504
rect 5686 17448 5691 17504
rect 0 17446 5691 17448
rect 0 17416 800 17446
rect 5625 17443 5691 17446
rect 10133 17506 10199 17509
rect 11789 17506 11855 17509
rect 13629 17506 13695 17509
rect 10133 17504 13695 17506
rect 10133 17448 10138 17504
rect 10194 17448 11794 17504
rect 11850 17448 13634 17504
rect 13690 17448 13695 17504
rect 10133 17446 13695 17448
rect 10133 17443 10199 17446
rect 11789 17443 11855 17446
rect 13629 17443 13695 17446
rect 8210 17440 8526 17441
rect 8210 17376 8216 17440
rect 8280 17376 8296 17440
rect 8360 17376 8376 17440
rect 8440 17376 8456 17440
rect 8520 17376 8526 17440
rect 8210 17375 8526 17376
rect 16210 17440 16526 17441
rect 16210 17376 16216 17440
rect 16280 17376 16296 17440
rect 16360 17376 16376 17440
rect 16440 17376 16456 17440
rect 16520 17376 16526 17440
rect 16210 17375 16526 17376
rect 24210 17440 24526 17441
rect 24210 17376 24216 17440
rect 24280 17376 24296 17440
rect 24360 17376 24376 17440
rect 24440 17376 24456 17440
rect 24520 17376 24526 17440
rect 24210 17375 24526 17376
rect 9213 17370 9279 17373
rect 12709 17370 12775 17373
rect 9213 17368 12775 17370
rect 9213 17312 9218 17368
rect 9274 17312 12714 17368
rect 12770 17312 12775 17368
rect 9213 17310 12775 17312
rect 9213 17307 9279 17310
rect 12709 17307 12775 17310
rect 10225 17234 10291 17237
rect 10593 17234 10659 17237
rect 15377 17234 15443 17237
rect 10225 17232 15443 17234
rect 10225 17176 10230 17232
rect 10286 17176 10598 17232
rect 10654 17176 15382 17232
rect 15438 17176 15443 17232
rect 10225 17174 15443 17176
rect 10225 17171 10291 17174
rect 10593 17171 10659 17174
rect 15377 17171 15443 17174
rect 9857 17098 9923 17101
rect 13537 17098 13603 17101
rect 9857 17096 13603 17098
rect 9857 17040 9862 17096
rect 9918 17040 13542 17096
rect 13598 17040 13603 17096
rect 9857 17038 13603 17040
rect 9857 17035 9923 17038
rect 13537 17035 13603 17038
rect 12065 16962 12131 16965
rect 11654 16960 12131 16962
rect 11654 16904 12070 16960
rect 12126 16904 12131 16960
rect 11654 16902 12131 16904
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 11654 16829 11714 16902
rect 12065 16899 12131 16902
rect 12210 16896 12526 16897
rect 12210 16832 12216 16896
rect 12280 16832 12296 16896
rect 12360 16832 12376 16896
rect 12440 16832 12456 16896
rect 12520 16832 12526 16896
rect 12210 16831 12526 16832
rect 20210 16896 20526 16897
rect 20210 16832 20216 16896
rect 20280 16832 20296 16896
rect 20360 16832 20376 16896
rect 20440 16832 20456 16896
rect 20520 16832 20526 16896
rect 20210 16831 20526 16832
rect 11605 16824 11714 16829
rect 11605 16768 11610 16824
rect 11666 16768 11714 16824
rect 11605 16766 11714 16768
rect 11605 16763 11671 16766
rect 10409 16690 10475 16693
rect 12065 16690 12131 16693
rect 14457 16690 14523 16693
rect 10409 16688 14523 16690
rect 10409 16632 10414 16688
rect 10470 16632 12070 16688
rect 12126 16632 14462 16688
rect 14518 16632 14523 16688
rect 10409 16630 14523 16632
rect 10409 16627 10475 16630
rect 12065 16627 12131 16630
rect 14457 16627 14523 16630
rect 11237 16554 11303 16557
rect 12157 16554 12223 16557
rect 11237 16552 12223 16554
rect 11237 16496 11242 16552
rect 11298 16496 12162 16552
rect 12218 16496 12223 16552
rect 11237 16494 12223 16496
rect 11237 16491 11303 16494
rect 12157 16491 12223 16494
rect 0 16418 800 16448
rect 7373 16418 7439 16421
rect 0 16416 7439 16418
rect 0 16360 7378 16416
rect 7434 16360 7439 16416
rect 0 16358 7439 16360
rect 0 16328 800 16358
rect 7373 16355 7439 16358
rect 9765 16418 9831 16421
rect 11881 16418 11947 16421
rect 9765 16416 11947 16418
rect 9765 16360 9770 16416
rect 9826 16360 11886 16416
rect 11942 16360 11947 16416
rect 9765 16358 11947 16360
rect 9765 16355 9831 16358
rect 11881 16355 11947 16358
rect 8210 16352 8526 16353
rect 8210 16288 8216 16352
rect 8280 16288 8296 16352
rect 8360 16288 8376 16352
rect 8440 16288 8456 16352
rect 8520 16288 8526 16352
rect 8210 16287 8526 16288
rect 16210 16352 16526 16353
rect 16210 16288 16216 16352
rect 16280 16288 16296 16352
rect 16360 16288 16376 16352
rect 16440 16288 16456 16352
rect 16520 16288 16526 16352
rect 16210 16287 16526 16288
rect 24210 16352 24526 16353
rect 24210 16288 24216 16352
rect 24280 16288 24296 16352
rect 24360 16288 24376 16352
rect 24440 16288 24456 16352
rect 24520 16288 24526 16352
rect 24210 16287 24526 16288
rect 11605 16284 11671 16285
rect 11605 16282 11652 16284
rect 11560 16280 11652 16282
rect 11560 16224 11610 16280
rect 11560 16222 11652 16224
rect 11605 16220 11652 16222
rect 11716 16220 11722 16284
rect 11605 16219 11671 16220
rect 10961 16146 11027 16149
rect 17033 16146 17099 16149
rect 10961 16144 17099 16146
rect 10961 16088 10966 16144
rect 11022 16088 17038 16144
rect 17094 16088 17099 16144
rect 10961 16086 17099 16088
rect 10961 16083 11027 16086
rect 17033 16083 17099 16086
rect 24853 16146 24919 16149
rect 26200 16146 27000 16176
rect 24853 16144 27000 16146
rect 24853 16088 24858 16144
rect 24914 16088 27000 16144
rect 24853 16086 27000 16088
rect 24853 16083 24919 16086
rect 26200 16056 27000 16086
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 12210 15808 12526 15809
rect 12210 15744 12216 15808
rect 12280 15744 12296 15808
rect 12360 15744 12376 15808
rect 12440 15744 12456 15808
rect 12520 15744 12526 15808
rect 12210 15743 12526 15744
rect 20210 15808 20526 15809
rect 20210 15744 20216 15808
rect 20280 15744 20296 15808
rect 20360 15744 20376 15808
rect 20440 15744 20456 15808
rect 20520 15744 20526 15808
rect 20210 15743 20526 15744
rect 0 15330 800 15360
rect 6913 15330 6979 15333
rect 0 15328 6979 15330
rect 0 15272 6918 15328
rect 6974 15272 6979 15328
rect 0 15270 6979 15272
rect 0 15240 800 15270
rect 6913 15267 6979 15270
rect 8210 15264 8526 15265
rect 8210 15200 8216 15264
rect 8280 15200 8296 15264
rect 8360 15200 8376 15264
rect 8440 15200 8456 15264
rect 8520 15200 8526 15264
rect 8210 15199 8526 15200
rect 16210 15264 16526 15265
rect 16210 15200 16216 15264
rect 16280 15200 16296 15264
rect 16360 15200 16376 15264
rect 16440 15200 16456 15264
rect 16520 15200 16526 15264
rect 16210 15199 16526 15200
rect 24210 15264 24526 15265
rect 24210 15200 24216 15264
rect 24280 15200 24296 15264
rect 24360 15200 24376 15264
rect 24440 15200 24456 15264
rect 24520 15200 24526 15264
rect 24210 15199 24526 15200
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 12210 14720 12526 14721
rect 12210 14656 12216 14720
rect 12280 14656 12296 14720
rect 12360 14656 12376 14720
rect 12440 14656 12456 14720
rect 12520 14656 12526 14720
rect 12210 14655 12526 14656
rect 20210 14720 20526 14721
rect 20210 14656 20216 14720
rect 20280 14656 20296 14720
rect 20360 14656 20376 14720
rect 20440 14656 20456 14720
rect 20520 14656 20526 14720
rect 20210 14655 20526 14656
rect 0 14242 800 14272
rect 6453 14242 6519 14245
rect 0 14240 6519 14242
rect 0 14184 6458 14240
rect 6514 14184 6519 14240
rect 0 14182 6519 14184
rect 0 14152 800 14182
rect 6453 14179 6519 14182
rect 8210 14176 8526 14177
rect 8210 14112 8216 14176
rect 8280 14112 8296 14176
rect 8360 14112 8376 14176
rect 8440 14112 8456 14176
rect 8520 14112 8526 14176
rect 8210 14111 8526 14112
rect 16210 14176 16526 14177
rect 16210 14112 16216 14176
rect 16280 14112 16296 14176
rect 16360 14112 16376 14176
rect 16440 14112 16456 14176
rect 16520 14112 16526 14176
rect 16210 14111 16526 14112
rect 24210 14176 24526 14177
rect 24210 14112 24216 14176
rect 24280 14112 24296 14176
rect 24360 14112 24376 14176
rect 24440 14112 24456 14176
rect 24520 14112 24526 14176
rect 24210 14111 24526 14112
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 12210 13632 12526 13633
rect 12210 13568 12216 13632
rect 12280 13568 12296 13632
rect 12360 13568 12376 13632
rect 12440 13568 12456 13632
rect 12520 13568 12526 13632
rect 12210 13567 12526 13568
rect 20210 13632 20526 13633
rect 20210 13568 20216 13632
rect 20280 13568 20296 13632
rect 20360 13568 20376 13632
rect 20440 13568 20456 13632
rect 20520 13568 20526 13632
rect 20210 13567 20526 13568
rect 0 13154 800 13184
rect 0 13094 2790 13154
rect 0 13064 800 13094
rect 2730 12882 2790 13094
rect 8210 13088 8526 13089
rect 8210 13024 8216 13088
rect 8280 13024 8296 13088
rect 8360 13024 8376 13088
rect 8440 13024 8456 13088
rect 8520 13024 8526 13088
rect 8210 13023 8526 13024
rect 16210 13088 16526 13089
rect 16210 13024 16216 13088
rect 16280 13024 16296 13088
rect 16360 13024 16376 13088
rect 16440 13024 16456 13088
rect 16520 13024 16526 13088
rect 16210 13023 16526 13024
rect 24210 13088 24526 13089
rect 24210 13024 24216 13088
rect 24280 13024 24296 13088
rect 24360 13024 24376 13088
rect 24440 13024 24456 13088
rect 24520 13024 24526 13088
rect 24210 13023 24526 13024
rect 13629 12882 13695 12885
rect 2730 12880 13695 12882
rect 2730 12824 13634 12880
rect 13690 12824 13695 12880
rect 2730 12822 13695 12824
rect 13629 12819 13695 12822
rect 24945 12610 25011 12613
rect 26200 12610 27000 12640
rect 24945 12608 27000 12610
rect 24945 12552 24950 12608
rect 25006 12552 27000 12608
rect 24945 12550 27000 12552
rect 24945 12547 25011 12550
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 12210 12544 12526 12545
rect 12210 12480 12216 12544
rect 12280 12480 12296 12544
rect 12360 12480 12376 12544
rect 12440 12480 12456 12544
rect 12520 12480 12526 12544
rect 12210 12479 12526 12480
rect 20210 12544 20526 12545
rect 20210 12480 20216 12544
rect 20280 12480 20296 12544
rect 20360 12480 20376 12544
rect 20440 12480 20456 12544
rect 20520 12480 20526 12544
rect 26200 12520 27000 12550
rect 20210 12479 20526 12480
rect 10685 12202 10751 12205
rect 2730 12200 10751 12202
rect 2730 12144 10690 12200
rect 10746 12144 10751 12200
rect 2730 12142 10751 12144
rect 0 12066 800 12096
rect 2730 12066 2790 12142
rect 10685 12139 10751 12142
rect 0 12006 2790 12066
rect 0 11976 800 12006
rect 8210 12000 8526 12001
rect 8210 11936 8216 12000
rect 8280 11936 8296 12000
rect 8360 11936 8376 12000
rect 8440 11936 8456 12000
rect 8520 11936 8526 12000
rect 8210 11935 8526 11936
rect 16210 12000 16526 12001
rect 16210 11936 16216 12000
rect 16280 11936 16296 12000
rect 16360 11936 16376 12000
rect 16440 11936 16456 12000
rect 16520 11936 16526 12000
rect 16210 11935 16526 11936
rect 24210 12000 24526 12001
rect 24210 11936 24216 12000
rect 24280 11936 24296 12000
rect 24360 11936 24376 12000
rect 24440 11936 24456 12000
rect 24520 11936 24526 12000
rect 24210 11935 24526 11936
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 12210 11456 12526 11457
rect 12210 11392 12216 11456
rect 12280 11392 12296 11456
rect 12360 11392 12376 11456
rect 12440 11392 12456 11456
rect 12520 11392 12526 11456
rect 12210 11391 12526 11392
rect 20210 11456 20526 11457
rect 20210 11392 20216 11456
rect 20280 11392 20296 11456
rect 20360 11392 20376 11456
rect 20440 11392 20456 11456
rect 20520 11392 20526 11456
rect 20210 11391 20526 11392
rect 0 10978 800 11008
rect 1301 10978 1367 10981
rect 0 10976 1367 10978
rect 0 10920 1306 10976
rect 1362 10920 1367 10976
rect 0 10918 1367 10920
rect 0 10888 800 10918
rect 1301 10915 1367 10918
rect 8210 10912 8526 10913
rect 8210 10848 8216 10912
rect 8280 10848 8296 10912
rect 8360 10848 8376 10912
rect 8440 10848 8456 10912
rect 8520 10848 8526 10912
rect 8210 10847 8526 10848
rect 16210 10912 16526 10913
rect 16210 10848 16216 10912
rect 16280 10848 16296 10912
rect 16360 10848 16376 10912
rect 16440 10848 16456 10912
rect 16520 10848 16526 10912
rect 16210 10847 16526 10848
rect 24210 10912 24526 10913
rect 24210 10848 24216 10912
rect 24280 10848 24296 10912
rect 24360 10848 24376 10912
rect 24440 10848 24456 10912
rect 24520 10848 24526 10912
rect 24210 10847 24526 10848
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 12210 10368 12526 10369
rect 12210 10304 12216 10368
rect 12280 10304 12296 10368
rect 12360 10304 12376 10368
rect 12440 10304 12456 10368
rect 12520 10304 12526 10368
rect 12210 10303 12526 10304
rect 20210 10368 20526 10369
rect 20210 10304 20216 10368
rect 20280 10304 20296 10368
rect 20360 10304 20376 10368
rect 20440 10304 20456 10368
rect 20520 10304 20526 10368
rect 20210 10303 20526 10304
rect 0 9890 800 9920
rect 6177 9890 6243 9893
rect 0 9888 6243 9890
rect 0 9832 6182 9888
rect 6238 9832 6243 9888
rect 0 9830 6243 9832
rect 0 9800 800 9830
rect 6177 9827 6243 9830
rect 8210 9824 8526 9825
rect 8210 9760 8216 9824
rect 8280 9760 8296 9824
rect 8360 9760 8376 9824
rect 8440 9760 8456 9824
rect 8520 9760 8526 9824
rect 8210 9759 8526 9760
rect 16210 9824 16526 9825
rect 16210 9760 16216 9824
rect 16280 9760 16296 9824
rect 16360 9760 16376 9824
rect 16440 9760 16456 9824
rect 16520 9760 16526 9824
rect 16210 9759 16526 9760
rect 24210 9824 24526 9825
rect 24210 9760 24216 9824
rect 24280 9760 24296 9824
rect 24360 9760 24376 9824
rect 24440 9760 24456 9824
rect 24520 9760 24526 9824
rect 24210 9759 24526 9760
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 12210 9280 12526 9281
rect 12210 9216 12216 9280
rect 12280 9216 12296 9280
rect 12360 9216 12376 9280
rect 12440 9216 12456 9280
rect 12520 9216 12526 9280
rect 12210 9215 12526 9216
rect 20210 9280 20526 9281
rect 20210 9216 20216 9280
rect 20280 9216 20296 9280
rect 20360 9216 20376 9280
rect 20440 9216 20456 9280
rect 20520 9216 20526 9280
rect 20210 9215 20526 9216
rect 15929 9074 15995 9077
rect 26200 9074 27000 9104
rect 15929 9072 27000 9074
rect 15929 9016 15934 9072
rect 15990 9016 27000 9072
rect 15929 9014 27000 9016
rect 15929 9011 15995 9014
rect 26200 8984 27000 9014
rect 0 8802 800 8832
rect 1301 8802 1367 8805
rect 0 8800 1367 8802
rect 0 8744 1306 8800
rect 1362 8744 1367 8800
rect 0 8742 1367 8744
rect 0 8712 800 8742
rect 1301 8739 1367 8742
rect 8210 8736 8526 8737
rect 8210 8672 8216 8736
rect 8280 8672 8296 8736
rect 8360 8672 8376 8736
rect 8440 8672 8456 8736
rect 8520 8672 8526 8736
rect 8210 8671 8526 8672
rect 16210 8736 16526 8737
rect 16210 8672 16216 8736
rect 16280 8672 16296 8736
rect 16360 8672 16376 8736
rect 16440 8672 16456 8736
rect 16520 8672 16526 8736
rect 16210 8671 16526 8672
rect 24210 8736 24526 8737
rect 24210 8672 24216 8736
rect 24280 8672 24296 8736
rect 24360 8672 24376 8736
rect 24440 8672 24456 8736
rect 24520 8672 24526 8736
rect 24210 8671 24526 8672
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 12210 8192 12526 8193
rect 12210 8128 12216 8192
rect 12280 8128 12296 8192
rect 12360 8128 12376 8192
rect 12440 8128 12456 8192
rect 12520 8128 12526 8192
rect 12210 8127 12526 8128
rect 20210 8192 20526 8193
rect 20210 8128 20216 8192
rect 20280 8128 20296 8192
rect 20360 8128 20376 8192
rect 20440 8128 20456 8192
rect 20520 8128 20526 8192
rect 20210 8127 20526 8128
rect 0 7714 800 7744
rect 4981 7714 5047 7717
rect 0 7712 5047 7714
rect 0 7656 4986 7712
rect 5042 7656 5047 7712
rect 0 7654 5047 7656
rect 0 7624 800 7654
rect 4981 7651 5047 7654
rect 8210 7648 8526 7649
rect 8210 7584 8216 7648
rect 8280 7584 8296 7648
rect 8360 7584 8376 7648
rect 8440 7584 8456 7648
rect 8520 7584 8526 7648
rect 8210 7583 8526 7584
rect 16210 7648 16526 7649
rect 16210 7584 16216 7648
rect 16280 7584 16296 7648
rect 16360 7584 16376 7648
rect 16440 7584 16456 7648
rect 16520 7584 16526 7648
rect 16210 7583 16526 7584
rect 24210 7648 24526 7649
rect 24210 7584 24216 7648
rect 24280 7584 24296 7648
rect 24360 7584 24376 7648
rect 24440 7584 24456 7648
rect 24520 7584 24526 7648
rect 24210 7583 24526 7584
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 12210 7104 12526 7105
rect 12210 7040 12216 7104
rect 12280 7040 12296 7104
rect 12360 7040 12376 7104
rect 12440 7040 12456 7104
rect 12520 7040 12526 7104
rect 12210 7039 12526 7040
rect 20210 7104 20526 7105
rect 20210 7040 20216 7104
rect 20280 7040 20296 7104
rect 20360 7040 20376 7104
rect 20440 7040 20456 7104
rect 20520 7040 20526 7104
rect 20210 7039 20526 7040
rect 0 6626 800 6656
rect 3325 6626 3391 6629
rect 0 6624 3391 6626
rect 0 6568 3330 6624
rect 3386 6568 3391 6624
rect 0 6566 3391 6568
rect 0 6536 800 6566
rect 3325 6563 3391 6566
rect 8210 6560 8526 6561
rect 8210 6496 8216 6560
rect 8280 6496 8296 6560
rect 8360 6496 8376 6560
rect 8440 6496 8456 6560
rect 8520 6496 8526 6560
rect 8210 6495 8526 6496
rect 16210 6560 16526 6561
rect 16210 6496 16216 6560
rect 16280 6496 16296 6560
rect 16360 6496 16376 6560
rect 16440 6496 16456 6560
rect 16520 6496 16526 6560
rect 16210 6495 16526 6496
rect 24210 6560 24526 6561
rect 24210 6496 24216 6560
rect 24280 6496 24296 6560
rect 24360 6496 24376 6560
rect 24440 6496 24456 6560
rect 24520 6496 24526 6560
rect 24210 6495 24526 6496
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 12210 6016 12526 6017
rect 12210 5952 12216 6016
rect 12280 5952 12296 6016
rect 12360 5952 12376 6016
rect 12440 5952 12456 6016
rect 12520 5952 12526 6016
rect 12210 5951 12526 5952
rect 20210 6016 20526 6017
rect 20210 5952 20216 6016
rect 20280 5952 20296 6016
rect 20360 5952 20376 6016
rect 20440 5952 20456 6016
rect 20520 5952 20526 6016
rect 20210 5951 20526 5952
rect 11421 5674 11487 5677
rect 15745 5674 15811 5677
rect 11421 5672 15811 5674
rect 11421 5616 11426 5672
rect 11482 5616 15750 5672
rect 15806 5616 15811 5672
rect 11421 5614 15811 5616
rect 11421 5611 11487 5614
rect 15745 5611 15811 5614
rect 0 5538 800 5568
rect 26200 5541 27000 5568
rect 3049 5538 3115 5541
rect 0 5536 3115 5538
rect 0 5480 3054 5536
rect 3110 5480 3115 5536
rect 0 5478 3115 5480
rect 0 5448 800 5478
rect 3049 5475 3115 5478
rect 26141 5536 27000 5541
rect 26141 5480 26146 5536
rect 26202 5480 27000 5536
rect 26141 5475 27000 5480
rect 8210 5472 8526 5473
rect 8210 5408 8216 5472
rect 8280 5408 8296 5472
rect 8360 5408 8376 5472
rect 8440 5408 8456 5472
rect 8520 5408 8526 5472
rect 8210 5407 8526 5408
rect 16210 5472 16526 5473
rect 16210 5408 16216 5472
rect 16280 5408 16296 5472
rect 16360 5408 16376 5472
rect 16440 5408 16456 5472
rect 16520 5408 16526 5472
rect 16210 5407 16526 5408
rect 24210 5472 24526 5473
rect 24210 5408 24216 5472
rect 24280 5408 24296 5472
rect 24360 5408 24376 5472
rect 24440 5408 24456 5472
rect 24520 5408 24526 5472
rect 26200 5448 27000 5475
rect 24210 5407 24526 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 12210 4928 12526 4929
rect 12210 4864 12216 4928
rect 12280 4864 12296 4928
rect 12360 4864 12376 4928
rect 12440 4864 12456 4928
rect 12520 4864 12526 4928
rect 12210 4863 12526 4864
rect 20210 4928 20526 4929
rect 20210 4864 20216 4928
rect 20280 4864 20296 4928
rect 20360 4864 20376 4928
rect 20440 4864 20456 4928
rect 20520 4864 20526 4928
rect 20210 4863 20526 4864
rect 0 4450 800 4480
rect 5073 4450 5139 4453
rect 0 4448 5139 4450
rect 0 4392 5078 4448
rect 5134 4392 5139 4448
rect 0 4390 5139 4392
rect 0 4360 800 4390
rect 5073 4387 5139 4390
rect 8210 4384 8526 4385
rect 8210 4320 8216 4384
rect 8280 4320 8296 4384
rect 8360 4320 8376 4384
rect 8440 4320 8456 4384
rect 8520 4320 8526 4384
rect 8210 4319 8526 4320
rect 16210 4384 16526 4385
rect 16210 4320 16216 4384
rect 16280 4320 16296 4384
rect 16360 4320 16376 4384
rect 16440 4320 16456 4384
rect 16520 4320 16526 4384
rect 16210 4319 16526 4320
rect 24210 4384 24526 4385
rect 24210 4320 24216 4384
rect 24280 4320 24296 4384
rect 24360 4320 24376 4384
rect 24440 4320 24456 4384
rect 24520 4320 24526 4384
rect 24210 4319 24526 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 12210 3840 12526 3841
rect 12210 3776 12216 3840
rect 12280 3776 12296 3840
rect 12360 3776 12376 3840
rect 12440 3776 12456 3840
rect 12520 3776 12526 3840
rect 12210 3775 12526 3776
rect 20210 3840 20526 3841
rect 20210 3776 20216 3840
rect 20280 3776 20296 3840
rect 20360 3776 20376 3840
rect 20440 3776 20456 3840
rect 20520 3776 20526 3840
rect 20210 3775 20526 3776
rect 0 3362 800 3392
rect 5901 3362 5967 3365
rect 0 3360 5967 3362
rect 0 3304 5906 3360
rect 5962 3304 5967 3360
rect 0 3302 5967 3304
rect 0 3272 800 3302
rect 5901 3299 5967 3302
rect 8210 3296 8526 3297
rect 8210 3232 8216 3296
rect 8280 3232 8296 3296
rect 8360 3232 8376 3296
rect 8440 3232 8456 3296
rect 8520 3232 8526 3296
rect 8210 3231 8526 3232
rect 16210 3296 16526 3297
rect 16210 3232 16216 3296
rect 16280 3232 16296 3296
rect 16360 3232 16376 3296
rect 16440 3232 16456 3296
rect 16520 3232 16526 3296
rect 16210 3231 16526 3232
rect 24210 3296 24526 3297
rect 24210 3232 24216 3296
rect 24280 3232 24296 3296
rect 24360 3232 24376 3296
rect 24440 3232 24456 3296
rect 24520 3232 24526 3296
rect 24210 3231 24526 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 12210 2752 12526 2753
rect 12210 2688 12216 2752
rect 12280 2688 12296 2752
rect 12360 2688 12376 2752
rect 12440 2688 12456 2752
rect 12520 2688 12526 2752
rect 12210 2687 12526 2688
rect 20210 2752 20526 2753
rect 20210 2688 20216 2752
rect 20280 2688 20296 2752
rect 20360 2688 20376 2752
rect 20440 2688 20456 2752
rect 20520 2688 20526 2752
rect 20210 2687 20526 2688
rect 197 2546 263 2549
rect 197 2544 1042 2546
rect 197 2488 202 2544
rect 258 2488 1042 2544
rect 197 2486 1042 2488
rect 197 2483 263 2486
rect 0 2274 800 2304
rect 982 2274 1042 2486
rect 0 2214 1042 2274
rect 0 2184 800 2214
rect 8210 2208 8526 2209
rect 8210 2144 8216 2208
rect 8280 2144 8296 2208
rect 8360 2144 8376 2208
rect 8440 2144 8456 2208
rect 8520 2144 8526 2208
rect 8210 2143 8526 2144
rect 16210 2208 16526 2209
rect 16210 2144 16216 2208
rect 16280 2144 16296 2208
rect 16360 2144 16376 2208
rect 16440 2144 16456 2208
rect 16520 2144 16526 2208
rect 16210 2143 16526 2144
rect 24210 2208 24526 2209
rect 24210 2144 24216 2208
rect 24280 2144 24296 2208
rect 24360 2144 24376 2208
rect 24440 2144 24456 2208
rect 24520 2144 24526 2208
rect 24210 2143 24526 2144
rect 26200 2005 27000 2032
rect 26141 2000 27000 2005
rect 26141 1944 26146 2000
rect 26202 1944 27000 2000
rect 26141 1939 27000 1944
rect 26200 1912 27000 1939
rect 4210 1664 4526 1665
rect 4210 1600 4216 1664
rect 4280 1600 4296 1664
rect 4360 1600 4376 1664
rect 4440 1600 4456 1664
rect 4520 1600 4526 1664
rect 4210 1599 4526 1600
rect 12210 1664 12526 1665
rect 12210 1600 12216 1664
rect 12280 1600 12296 1664
rect 12360 1600 12376 1664
rect 12440 1600 12456 1664
rect 12520 1600 12526 1664
rect 12210 1599 12526 1600
rect 20210 1664 20526 1665
rect 20210 1600 20216 1664
rect 20280 1600 20296 1664
rect 20360 1600 20376 1664
rect 20440 1600 20456 1664
rect 20520 1600 20526 1664
rect 20210 1599 20526 1600
rect 841 1322 907 1325
rect 798 1320 907 1322
rect 798 1264 846 1320
rect 902 1264 907 1320
rect 798 1259 907 1264
rect 798 1216 858 1259
rect 0 1126 858 1216
rect 0 1096 800 1126
rect 8210 1120 8526 1121
rect 8210 1056 8216 1120
rect 8280 1056 8296 1120
rect 8360 1056 8376 1120
rect 8440 1056 8456 1120
rect 8520 1056 8526 1120
rect 8210 1055 8526 1056
rect 16210 1120 16526 1121
rect 16210 1056 16216 1120
rect 16280 1056 16296 1120
rect 16360 1056 16376 1120
rect 16440 1056 16456 1120
rect 16520 1056 16526 1120
rect 16210 1055 16526 1056
rect 24210 1120 24526 1121
rect 24210 1056 24216 1120
rect 24280 1056 24296 1120
rect 24360 1056 24376 1120
rect 24440 1056 24456 1120
rect 24520 1056 24526 1120
rect 24210 1055 24526 1056
<< via3 >>
rect 8216 20700 8280 20704
rect 8216 20644 8220 20700
rect 8220 20644 8276 20700
rect 8276 20644 8280 20700
rect 8216 20640 8280 20644
rect 8296 20700 8360 20704
rect 8296 20644 8300 20700
rect 8300 20644 8356 20700
rect 8356 20644 8360 20700
rect 8296 20640 8360 20644
rect 8376 20700 8440 20704
rect 8376 20644 8380 20700
rect 8380 20644 8436 20700
rect 8436 20644 8440 20700
rect 8376 20640 8440 20644
rect 8456 20700 8520 20704
rect 8456 20644 8460 20700
rect 8460 20644 8516 20700
rect 8516 20644 8520 20700
rect 8456 20640 8520 20644
rect 16216 20700 16280 20704
rect 16216 20644 16220 20700
rect 16220 20644 16276 20700
rect 16276 20644 16280 20700
rect 16216 20640 16280 20644
rect 16296 20700 16360 20704
rect 16296 20644 16300 20700
rect 16300 20644 16356 20700
rect 16356 20644 16360 20700
rect 16296 20640 16360 20644
rect 16376 20700 16440 20704
rect 16376 20644 16380 20700
rect 16380 20644 16436 20700
rect 16436 20644 16440 20700
rect 16376 20640 16440 20644
rect 16456 20700 16520 20704
rect 16456 20644 16460 20700
rect 16460 20644 16516 20700
rect 16516 20644 16520 20700
rect 16456 20640 16520 20644
rect 24216 20700 24280 20704
rect 24216 20644 24220 20700
rect 24220 20644 24276 20700
rect 24276 20644 24280 20700
rect 24216 20640 24280 20644
rect 24296 20700 24360 20704
rect 24296 20644 24300 20700
rect 24300 20644 24356 20700
rect 24356 20644 24360 20700
rect 24296 20640 24360 20644
rect 24376 20700 24440 20704
rect 24376 20644 24380 20700
rect 24380 20644 24436 20700
rect 24436 20644 24440 20700
rect 24376 20640 24440 20644
rect 24456 20700 24520 20704
rect 24456 20644 24460 20700
rect 24460 20644 24516 20700
rect 24516 20644 24520 20700
rect 24456 20640 24520 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 12216 20156 12280 20160
rect 12216 20100 12220 20156
rect 12220 20100 12276 20156
rect 12276 20100 12280 20156
rect 12216 20096 12280 20100
rect 12296 20156 12360 20160
rect 12296 20100 12300 20156
rect 12300 20100 12356 20156
rect 12356 20100 12360 20156
rect 12296 20096 12360 20100
rect 12376 20156 12440 20160
rect 12376 20100 12380 20156
rect 12380 20100 12436 20156
rect 12436 20100 12440 20156
rect 12376 20096 12440 20100
rect 12456 20156 12520 20160
rect 12456 20100 12460 20156
rect 12460 20100 12516 20156
rect 12516 20100 12520 20156
rect 12456 20096 12520 20100
rect 20216 20156 20280 20160
rect 20216 20100 20220 20156
rect 20220 20100 20276 20156
rect 20276 20100 20280 20156
rect 20216 20096 20280 20100
rect 20296 20156 20360 20160
rect 20296 20100 20300 20156
rect 20300 20100 20356 20156
rect 20356 20100 20360 20156
rect 20296 20096 20360 20100
rect 20376 20156 20440 20160
rect 20376 20100 20380 20156
rect 20380 20100 20436 20156
rect 20436 20100 20440 20156
rect 20376 20096 20440 20100
rect 20456 20156 20520 20160
rect 20456 20100 20460 20156
rect 20460 20100 20516 20156
rect 20516 20100 20520 20156
rect 20456 20096 20520 20100
rect 8216 19612 8280 19616
rect 8216 19556 8220 19612
rect 8220 19556 8276 19612
rect 8276 19556 8280 19612
rect 8216 19552 8280 19556
rect 8296 19612 8360 19616
rect 8296 19556 8300 19612
rect 8300 19556 8356 19612
rect 8356 19556 8360 19612
rect 8296 19552 8360 19556
rect 8376 19612 8440 19616
rect 8376 19556 8380 19612
rect 8380 19556 8436 19612
rect 8436 19556 8440 19612
rect 8376 19552 8440 19556
rect 8456 19612 8520 19616
rect 8456 19556 8460 19612
rect 8460 19556 8516 19612
rect 8516 19556 8520 19612
rect 8456 19552 8520 19556
rect 16216 19612 16280 19616
rect 16216 19556 16220 19612
rect 16220 19556 16276 19612
rect 16276 19556 16280 19612
rect 16216 19552 16280 19556
rect 16296 19612 16360 19616
rect 16296 19556 16300 19612
rect 16300 19556 16356 19612
rect 16356 19556 16360 19612
rect 16296 19552 16360 19556
rect 16376 19612 16440 19616
rect 16376 19556 16380 19612
rect 16380 19556 16436 19612
rect 16436 19556 16440 19612
rect 16376 19552 16440 19556
rect 16456 19612 16520 19616
rect 16456 19556 16460 19612
rect 16460 19556 16516 19612
rect 16516 19556 16520 19612
rect 16456 19552 16520 19556
rect 24216 19612 24280 19616
rect 24216 19556 24220 19612
rect 24220 19556 24276 19612
rect 24276 19556 24280 19612
rect 24216 19552 24280 19556
rect 24296 19612 24360 19616
rect 24296 19556 24300 19612
rect 24300 19556 24356 19612
rect 24356 19556 24360 19612
rect 24296 19552 24360 19556
rect 24376 19612 24440 19616
rect 24376 19556 24380 19612
rect 24380 19556 24436 19612
rect 24436 19556 24440 19612
rect 24376 19552 24440 19556
rect 24456 19612 24520 19616
rect 24456 19556 24460 19612
rect 24460 19556 24516 19612
rect 24516 19556 24520 19612
rect 24456 19552 24520 19556
rect 11468 19076 11532 19140
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 12216 19068 12280 19072
rect 12216 19012 12220 19068
rect 12220 19012 12276 19068
rect 12276 19012 12280 19068
rect 12216 19008 12280 19012
rect 12296 19068 12360 19072
rect 12296 19012 12300 19068
rect 12300 19012 12356 19068
rect 12356 19012 12360 19068
rect 12296 19008 12360 19012
rect 12376 19068 12440 19072
rect 12376 19012 12380 19068
rect 12380 19012 12436 19068
rect 12436 19012 12440 19068
rect 12376 19008 12440 19012
rect 12456 19068 12520 19072
rect 12456 19012 12460 19068
rect 12460 19012 12516 19068
rect 12516 19012 12520 19068
rect 12456 19008 12520 19012
rect 20216 19068 20280 19072
rect 20216 19012 20220 19068
rect 20220 19012 20276 19068
rect 20276 19012 20280 19068
rect 20216 19008 20280 19012
rect 20296 19068 20360 19072
rect 20296 19012 20300 19068
rect 20300 19012 20356 19068
rect 20356 19012 20360 19068
rect 20296 19008 20360 19012
rect 20376 19068 20440 19072
rect 20376 19012 20380 19068
rect 20380 19012 20436 19068
rect 20436 19012 20440 19068
rect 20376 19008 20440 19012
rect 20456 19068 20520 19072
rect 20456 19012 20460 19068
rect 20460 19012 20516 19068
rect 20516 19012 20520 19068
rect 20456 19008 20520 19012
rect 11652 18864 11716 18868
rect 11652 18808 11702 18864
rect 11702 18808 11716 18864
rect 11652 18804 11716 18808
rect 8216 18524 8280 18528
rect 8216 18468 8220 18524
rect 8220 18468 8276 18524
rect 8276 18468 8280 18524
rect 8216 18464 8280 18468
rect 8296 18524 8360 18528
rect 8296 18468 8300 18524
rect 8300 18468 8356 18524
rect 8356 18468 8360 18524
rect 8296 18464 8360 18468
rect 8376 18524 8440 18528
rect 8376 18468 8380 18524
rect 8380 18468 8436 18524
rect 8436 18468 8440 18524
rect 8376 18464 8440 18468
rect 8456 18524 8520 18528
rect 8456 18468 8460 18524
rect 8460 18468 8516 18524
rect 8516 18468 8520 18524
rect 8456 18464 8520 18468
rect 16216 18524 16280 18528
rect 16216 18468 16220 18524
rect 16220 18468 16276 18524
rect 16276 18468 16280 18524
rect 16216 18464 16280 18468
rect 16296 18524 16360 18528
rect 16296 18468 16300 18524
rect 16300 18468 16356 18524
rect 16356 18468 16360 18524
rect 16296 18464 16360 18468
rect 16376 18524 16440 18528
rect 16376 18468 16380 18524
rect 16380 18468 16436 18524
rect 16436 18468 16440 18524
rect 16376 18464 16440 18468
rect 16456 18524 16520 18528
rect 16456 18468 16460 18524
rect 16460 18468 16516 18524
rect 16516 18468 16520 18524
rect 16456 18464 16520 18468
rect 24216 18524 24280 18528
rect 24216 18468 24220 18524
rect 24220 18468 24276 18524
rect 24276 18468 24280 18524
rect 24216 18464 24280 18468
rect 24296 18524 24360 18528
rect 24296 18468 24300 18524
rect 24300 18468 24356 18524
rect 24356 18468 24360 18524
rect 24296 18464 24360 18468
rect 24376 18524 24440 18528
rect 24376 18468 24380 18524
rect 24380 18468 24436 18524
rect 24436 18468 24440 18524
rect 24376 18464 24440 18468
rect 24456 18524 24520 18528
rect 24456 18468 24460 18524
rect 24460 18468 24516 18524
rect 24516 18468 24520 18524
rect 24456 18464 24520 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 12216 17980 12280 17984
rect 12216 17924 12220 17980
rect 12220 17924 12276 17980
rect 12276 17924 12280 17980
rect 12216 17920 12280 17924
rect 12296 17980 12360 17984
rect 12296 17924 12300 17980
rect 12300 17924 12356 17980
rect 12356 17924 12360 17980
rect 12296 17920 12360 17924
rect 12376 17980 12440 17984
rect 12376 17924 12380 17980
rect 12380 17924 12436 17980
rect 12436 17924 12440 17980
rect 12376 17920 12440 17924
rect 12456 17980 12520 17984
rect 12456 17924 12460 17980
rect 12460 17924 12516 17980
rect 12516 17924 12520 17980
rect 12456 17920 12520 17924
rect 20216 17980 20280 17984
rect 20216 17924 20220 17980
rect 20220 17924 20276 17980
rect 20276 17924 20280 17980
rect 20216 17920 20280 17924
rect 20296 17980 20360 17984
rect 20296 17924 20300 17980
rect 20300 17924 20356 17980
rect 20356 17924 20360 17980
rect 20296 17920 20360 17924
rect 20376 17980 20440 17984
rect 20376 17924 20380 17980
rect 20380 17924 20436 17980
rect 20436 17924 20440 17980
rect 20376 17920 20440 17924
rect 20456 17980 20520 17984
rect 20456 17924 20460 17980
rect 20460 17924 20516 17980
rect 20516 17924 20520 17980
rect 20456 17920 20520 17924
rect 11468 17852 11532 17916
rect 8216 17436 8280 17440
rect 8216 17380 8220 17436
rect 8220 17380 8276 17436
rect 8276 17380 8280 17436
rect 8216 17376 8280 17380
rect 8296 17436 8360 17440
rect 8296 17380 8300 17436
rect 8300 17380 8356 17436
rect 8356 17380 8360 17436
rect 8296 17376 8360 17380
rect 8376 17436 8440 17440
rect 8376 17380 8380 17436
rect 8380 17380 8436 17436
rect 8436 17380 8440 17436
rect 8376 17376 8440 17380
rect 8456 17436 8520 17440
rect 8456 17380 8460 17436
rect 8460 17380 8516 17436
rect 8516 17380 8520 17436
rect 8456 17376 8520 17380
rect 16216 17436 16280 17440
rect 16216 17380 16220 17436
rect 16220 17380 16276 17436
rect 16276 17380 16280 17436
rect 16216 17376 16280 17380
rect 16296 17436 16360 17440
rect 16296 17380 16300 17436
rect 16300 17380 16356 17436
rect 16356 17380 16360 17436
rect 16296 17376 16360 17380
rect 16376 17436 16440 17440
rect 16376 17380 16380 17436
rect 16380 17380 16436 17436
rect 16436 17380 16440 17436
rect 16376 17376 16440 17380
rect 16456 17436 16520 17440
rect 16456 17380 16460 17436
rect 16460 17380 16516 17436
rect 16516 17380 16520 17436
rect 16456 17376 16520 17380
rect 24216 17436 24280 17440
rect 24216 17380 24220 17436
rect 24220 17380 24276 17436
rect 24276 17380 24280 17436
rect 24216 17376 24280 17380
rect 24296 17436 24360 17440
rect 24296 17380 24300 17436
rect 24300 17380 24356 17436
rect 24356 17380 24360 17436
rect 24296 17376 24360 17380
rect 24376 17436 24440 17440
rect 24376 17380 24380 17436
rect 24380 17380 24436 17436
rect 24436 17380 24440 17436
rect 24376 17376 24440 17380
rect 24456 17436 24520 17440
rect 24456 17380 24460 17436
rect 24460 17380 24516 17436
rect 24516 17380 24520 17436
rect 24456 17376 24520 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 12216 16892 12280 16896
rect 12216 16836 12220 16892
rect 12220 16836 12276 16892
rect 12276 16836 12280 16892
rect 12216 16832 12280 16836
rect 12296 16892 12360 16896
rect 12296 16836 12300 16892
rect 12300 16836 12356 16892
rect 12356 16836 12360 16892
rect 12296 16832 12360 16836
rect 12376 16892 12440 16896
rect 12376 16836 12380 16892
rect 12380 16836 12436 16892
rect 12436 16836 12440 16892
rect 12376 16832 12440 16836
rect 12456 16892 12520 16896
rect 12456 16836 12460 16892
rect 12460 16836 12516 16892
rect 12516 16836 12520 16892
rect 12456 16832 12520 16836
rect 20216 16892 20280 16896
rect 20216 16836 20220 16892
rect 20220 16836 20276 16892
rect 20276 16836 20280 16892
rect 20216 16832 20280 16836
rect 20296 16892 20360 16896
rect 20296 16836 20300 16892
rect 20300 16836 20356 16892
rect 20356 16836 20360 16892
rect 20296 16832 20360 16836
rect 20376 16892 20440 16896
rect 20376 16836 20380 16892
rect 20380 16836 20436 16892
rect 20436 16836 20440 16892
rect 20376 16832 20440 16836
rect 20456 16892 20520 16896
rect 20456 16836 20460 16892
rect 20460 16836 20516 16892
rect 20516 16836 20520 16892
rect 20456 16832 20520 16836
rect 8216 16348 8280 16352
rect 8216 16292 8220 16348
rect 8220 16292 8276 16348
rect 8276 16292 8280 16348
rect 8216 16288 8280 16292
rect 8296 16348 8360 16352
rect 8296 16292 8300 16348
rect 8300 16292 8356 16348
rect 8356 16292 8360 16348
rect 8296 16288 8360 16292
rect 8376 16348 8440 16352
rect 8376 16292 8380 16348
rect 8380 16292 8436 16348
rect 8436 16292 8440 16348
rect 8376 16288 8440 16292
rect 8456 16348 8520 16352
rect 8456 16292 8460 16348
rect 8460 16292 8516 16348
rect 8516 16292 8520 16348
rect 8456 16288 8520 16292
rect 16216 16348 16280 16352
rect 16216 16292 16220 16348
rect 16220 16292 16276 16348
rect 16276 16292 16280 16348
rect 16216 16288 16280 16292
rect 16296 16348 16360 16352
rect 16296 16292 16300 16348
rect 16300 16292 16356 16348
rect 16356 16292 16360 16348
rect 16296 16288 16360 16292
rect 16376 16348 16440 16352
rect 16376 16292 16380 16348
rect 16380 16292 16436 16348
rect 16436 16292 16440 16348
rect 16376 16288 16440 16292
rect 16456 16348 16520 16352
rect 16456 16292 16460 16348
rect 16460 16292 16516 16348
rect 16516 16292 16520 16348
rect 16456 16288 16520 16292
rect 24216 16348 24280 16352
rect 24216 16292 24220 16348
rect 24220 16292 24276 16348
rect 24276 16292 24280 16348
rect 24216 16288 24280 16292
rect 24296 16348 24360 16352
rect 24296 16292 24300 16348
rect 24300 16292 24356 16348
rect 24356 16292 24360 16348
rect 24296 16288 24360 16292
rect 24376 16348 24440 16352
rect 24376 16292 24380 16348
rect 24380 16292 24436 16348
rect 24436 16292 24440 16348
rect 24376 16288 24440 16292
rect 24456 16348 24520 16352
rect 24456 16292 24460 16348
rect 24460 16292 24516 16348
rect 24516 16292 24520 16348
rect 24456 16288 24520 16292
rect 11652 16280 11716 16284
rect 11652 16224 11666 16280
rect 11666 16224 11716 16280
rect 11652 16220 11716 16224
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 12216 15804 12280 15808
rect 12216 15748 12220 15804
rect 12220 15748 12276 15804
rect 12276 15748 12280 15804
rect 12216 15744 12280 15748
rect 12296 15804 12360 15808
rect 12296 15748 12300 15804
rect 12300 15748 12356 15804
rect 12356 15748 12360 15804
rect 12296 15744 12360 15748
rect 12376 15804 12440 15808
rect 12376 15748 12380 15804
rect 12380 15748 12436 15804
rect 12436 15748 12440 15804
rect 12376 15744 12440 15748
rect 12456 15804 12520 15808
rect 12456 15748 12460 15804
rect 12460 15748 12516 15804
rect 12516 15748 12520 15804
rect 12456 15744 12520 15748
rect 20216 15804 20280 15808
rect 20216 15748 20220 15804
rect 20220 15748 20276 15804
rect 20276 15748 20280 15804
rect 20216 15744 20280 15748
rect 20296 15804 20360 15808
rect 20296 15748 20300 15804
rect 20300 15748 20356 15804
rect 20356 15748 20360 15804
rect 20296 15744 20360 15748
rect 20376 15804 20440 15808
rect 20376 15748 20380 15804
rect 20380 15748 20436 15804
rect 20436 15748 20440 15804
rect 20376 15744 20440 15748
rect 20456 15804 20520 15808
rect 20456 15748 20460 15804
rect 20460 15748 20516 15804
rect 20516 15748 20520 15804
rect 20456 15744 20520 15748
rect 8216 15260 8280 15264
rect 8216 15204 8220 15260
rect 8220 15204 8276 15260
rect 8276 15204 8280 15260
rect 8216 15200 8280 15204
rect 8296 15260 8360 15264
rect 8296 15204 8300 15260
rect 8300 15204 8356 15260
rect 8356 15204 8360 15260
rect 8296 15200 8360 15204
rect 8376 15260 8440 15264
rect 8376 15204 8380 15260
rect 8380 15204 8436 15260
rect 8436 15204 8440 15260
rect 8376 15200 8440 15204
rect 8456 15260 8520 15264
rect 8456 15204 8460 15260
rect 8460 15204 8516 15260
rect 8516 15204 8520 15260
rect 8456 15200 8520 15204
rect 16216 15260 16280 15264
rect 16216 15204 16220 15260
rect 16220 15204 16276 15260
rect 16276 15204 16280 15260
rect 16216 15200 16280 15204
rect 16296 15260 16360 15264
rect 16296 15204 16300 15260
rect 16300 15204 16356 15260
rect 16356 15204 16360 15260
rect 16296 15200 16360 15204
rect 16376 15260 16440 15264
rect 16376 15204 16380 15260
rect 16380 15204 16436 15260
rect 16436 15204 16440 15260
rect 16376 15200 16440 15204
rect 16456 15260 16520 15264
rect 16456 15204 16460 15260
rect 16460 15204 16516 15260
rect 16516 15204 16520 15260
rect 16456 15200 16520 15204
rect 24216 15260 24280 15264
rect 24216 15204 24220 15260
rect 24220 15204 24276 15260
rect 24276 15204 24280 15260
rect 24216 15200 24280 15204
rect 24296 15260 24360 15264
rect 24296 15204 24300 15260
rect 24300 15204 24356 15260
rect 24356 15204 24360 15260
rect 24296 15200 24360 15204
rect 24376 15260 24440 15264
rect 24376 15204 24380 15260
rect 24380 15204 24436 15260
rect 24436 15204 24440 15260
rect 24376 15200 24440 15204
rect 24456 15260 24520 15264
rect 24456 15204 24460 15260
rect 24460 15204 24516 15260
rect 24516 15204 24520 15260
rect 24456 15200 24520 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 12216 14716 12280 14720
rect 12216 14660 12220 14716
rect 12220 14660 12276 14716
rect 12276 14660 12280 14716
rect 12216 14656 12280 14660
rect 12296 14716 12360 14720
rect 12296 14660 12300 14716
rect 12300 14660 12356 14716
rect 12356 14660 12360 14716
rect 12296 14656 12360 14660
rect 12376 14716 12440 14720
rect 12376 14660 12380 14716
rect 12380 14660 12436 14716
rect 12436 14660 12440 14716
rect 12376 14656 12440 14660
rect 12456 14716 12520 14720
rect 12456 14660 12460 14716
rect 12460 14660 12516 14716
rect 12516 14660 12520 14716
rect 12456 14656 12520 14660
rect 20216 14716 20280 14720
rect 20216 14660 20220 14716
rect 20220 14660 20276 14716
rect 20276 14660 20280 14716
rect 20216 14656 20280 14660
rect 20296 14716 20360 14720
rect 20296 14660 20300 14716
rect 20300 14660 20356 14716
rect 20356 14660 20360 14716
rect 20296 14656 20360 14660
rect 20376 14716 20440 14720
rect 20376 14660 20380 14716
rect 20380 14660 20436 14716
rect 20436 14660 20440 14716
rect 20376 14656 20440 14660
rect 20456 14716 20520 14720
rect 20456 14660 20460 14716
rect 20460 14660 20516 14716
rect 20516 14660 20520 14716
rect 20456 14656 20520 14660
rect 8216 14172 8280 14176
rect 8216 14116 8220 14172
rect 8220 14116 8276 14172
rect 8276 14116 8280 14172
rect 8216 14112 8280 14116
rect 8296 14172 8360 14176
rect 8296 14116 8300 14172
rect 8300 14116 8356 14172
rect 8356 14116 8360 14172
rect 8296 14112 8360 14116
rect 8376 14172 8440 14176
rect 8376 14116 8380 14172
rect 8380 14116 8436 14172
rect 8436 14116 8440 14172
rect 8376 14112 8440 14116
rect 8456 14172 8520 14176
rect 8456 14116 8460 14172
rect 8460 14116 8516 14172
rect 8516 14116 8520 14172
rect 8456 14112 8520 14116
rect 16216 14172 16280 14176
rect 16216 14116 16220 14172
rect 16220 14116 16276 14172
rect 16276 14116 16280 14172
rect 16216 14112 16280 14116
rect 16296 14172 16360 14176
rect 16296 14116 16300 14172
rect 16300 14116 16356 14172
rect 16356 14116 16360 14172
rect 16296 14112 16360 14116
rect 16376 14172 16440 14176
rect 16376 14116 16380 14172
rect 16380 14116 16436 14172
rect 16436 14116 16440 14172
rect 16376 14112 16440 14116
rect 16456 14172 16520 14176
rect 16456 14116 16460 14172
rect 16460 14116 16516 14172
rect 16516 14116 16520 14172
rect 16456 14112 16520 14116
rect 24216 14172 24280 14176
rect 24216 14116 24220 14172
rect 24220 14116 24276 14172
rect 24276 14116 24280 14172
rect 24216 14112 24280 14116
rect 24296 14172 24360 14176
rect 24296 14116 24300 14172
rect 24300 14116 24356 14172
rect 24356 14116 24360 14172
rect 24296 14112 24360 14116
rect 24376 14172 24440 14176
rect 24376 14116 24380 14172
rect 24380 14116 24436 14172
rect 24436 14116 24440 14172
rect 24376 14112 24440 14116
rect 24456 14172 24520 14176
rect 24456 14116 24460 14172
rect 24460 14116 24516 14172
rect 24516 14116 24520 14172
rect 24456 14112 24520 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 12216 13628 12280 13632
rect 12216 13572 12220 13628
rect 12220 13572 12276 13628
rect 12276 13572 12280 13628
rect 12216 13568 12280 13572
rect 12296 13628 12360 13632
rect 12296 13572 12300 13628
rect 12300 13572 12356 13628
rect 12356 13572 12360 13628
rect 12296 13568 12360 13572
rect 12376 13628 12440 13632
rect 12376 13572 12380 13628
rect 12380 13572 12436 13628
rect 12436 13572 12440 13628
rect 12376 13568 12440 13572
rect 12456 13628 12520 13632
rect 12456 13572 12460 13628
rect 12460 13572 12516 13628
rect 12516 13572 12520 13628
rect 12456 13568 12520 13572
rect 20216 13628 20280 13632
rect 20216 13572 20220 13628
rect 20220 13572 20276 13628
rect 20276 13572 20280 13628
rect 20216 13568 20280 13572
rect 20296 13628 20360 13632
rect 20296 13572 20300 13628
rect 20300 13572 20356 13628
rect 20356 13572 20360 13628
rect 20296 13568 20360 13572
rect 20376 13628 20440 13632
rect 20376 13572 20380 13628
rect 20380 13572 20436 13628
rect 20436 13572 20440 13628
rect 20376 13568 20440 13572
rect 20456 13628 20520 13632
rect 20456 13572 20460 13628
rect 20460 13572 20516 13628
rect 20516 13572 20520 13628
rect 20456 13568 20520 13572
rect 8216 13084 8280 13088
rect 8216 13028 8220 13084
rect 8220 13028 8276 13084
rect 8276 13028 8280 13084
rect 8216 13024 8280 13028
rect 8296 13084 8360 13088
rect 8296 13028 8300 13084
rect 8300 13028 8356 13084
rect 8356 13028 8360 13084
rect 8296 13024 8360 13028
rect 8376 13084 8440 13088
rect 8376 13028 8380 13084
rect 8380 13028 8436 13084
rect 8436 13028 8440 13084
rect 8376 13024 8440 13028
rect 8456 13084 8520 13088
rect 8456 13028 8460 13084
rect 8460 13028 8516 13084
rect 8516 13028 8520 13084
rect 8456 13024 8520 13028
rect 16216 13084 16280 13088
rect 16216 13028 16220 13084
rect 16220 13028 16276 13084
rect 16276 13028 16280 13084
rect 16216 13024 16280 13028
rect 16296 13084 16360 13088
rect 16296 13028 16300 13084
rect 16300 13028 16356 13084
rect 16356 13028 16360 13084
rect 16296 13024 16360 13028
rect 16376 13084 16440 13088
rect 16376 13028 16380 13084
rect 16380 13028 16436 13084
rect 16436 13028 16440 13084
rect 16376 13024 16440 13028
rect 16456 13084 16520 13088
rect 16456 13028 16460 13084
rect 16460 13028 16516 13084
rect 16516 13028 16520 13084
rect 16456 13024 16520 13028
rect 24216 13084 24280 13088
rect 24216 13028 24220 13084
rect 24220 13028 24276 13084
rect 24276 13028 24280 13084
rect 24216 13024 24280 13028
rect 24296 13084 24360 13088
rect 24296 13028 24300 13084
rect 24300 13028 24356 13084
rect 24356 13028 24360 13084
rect 24296 13024 24360 13028
rect 24376 13084 24440 13088
rect 24376 13028 24380 13084
rect 24380 13028 24436 13084
rect 24436 13028 24440 13084
rect 24376 13024 24440 13028
rect 24456 13084 24520 13088
rect 24456 13028 24460 13084
rect 24460 13028 24516 13084
rect 24516 13028 24520 13084
rect 24456 13024 24520 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 12216 12540 12280 12544
rect 12216 12484 12220 12540
rect 12220 12484 12276 12540
rect 12276 12484 12280 12540
rect 12216 12480 12280 12484
rect 12296 12540 12360 12544
rect 12296 12484 12300 12540
rect 12300 12484 12356 12540
rect 12356 12484 12360 12540
rect 12296 12480 12360 12484
rect 12376 12540 12440 12544
rect 12376 12484 12380 12540
rect 12380 12484 12436 12540
rect 12436 12484 12440 12540
rect 12376 12480 12440 12484
rect 12456 12540 12520 12544
rect 12456 12484 12460 12540
rect 12460 12484 12516 12540
rect 12516 12484 12520 12540
rect 12456 12480 12520 12484
rect 20216 12540 20280 12544
rect 20216 12484 20220 12540
rect 20220 12484 20276 12540
rect 20276 12484 20280 12540
rect 20216 12480 20280 12484
rect 20296 12540 20360 12544
rect 20296 12484 20300 12540
rect 20300 12484 20356 12540
rect 20356 12484 20360 12540
rect 20296 12480 20360 12484
rect 20376 12540 20440 12544
rect 20376 12484 20380 12540
rect 20380 12484 20436 12540
rect 20436 12484 20440 12540
rect 20376 12480 20440 12484
rect 20456 12540 20520 12544
rect 20456 12484 20460 12540
rect 20460 12484 20516 12540
rect 20516 12484 20520 12540
rect 20456 12480 20520 12484
rect 8216 11996 8280 12000
rect 8216 11940 8220 11996
rect 8220 11940 8276 11996
rect 8276 11940 8280 11996
rect 8216 11936 8280 11940
rect 8296 11996 8360 12000
rect 8296 11940 8300 11996
rect 8300 11940 8356 11996
rect 8356 11940 8360 11996
rect 8296 11936 8360 11940
rect 8376 11996 8440 12000
rect 8376 11940 8380 11996
rect 8380 11940 8436 11996
rect 8436 11940 8440 11996
rect 8376 11936 8440 11940
rect 8456 11996 8520 12000
rect 8456 11940 8460 11996
rect 8460 11940 8516 11996
rect 8516 11940 8520 11996
rect 8456 11936 8520 11940
rect 16216 11996 16280 12000
rect 16216 11940 16220 11996
rect 16220 11940 16276 11996
rect 16276 11940 16280 11996
rect 16216 11936 16280 11940
rect 16296 11996 16360 12000
rect 16296 11940 16300 11996
rect 16300 11940 16356 11996
rect 16356 11940 16360 11996
rect 16296 11936 16360 11940
rect 16376 11996 16440 12000
rect 16376 11940 16380 11996
rect 16380 11940 16436 11996
rect 16436 11940 16440 11996
rect 16376 11936 16440 11940
rect 16456 11996 16520 12000
rect 16456 11940 16460 11996
rect 16460 11940 16516 11996
rect 16516 11940 16520 11996
rect 16456 11936 16520 11940
rect 24216 11996 24280 12000
rect 24216 11940 24220 11996
rect 24220 11940 24276 11996
rect 24276 11940 24280 11996
rect 24216 11936 24280 11940
rect 24296 11996 24360 12000
rect 24296 11940 24300 11996
rect 24300 11940 24356 11996
rect 24356 11940 24360 11996
rect 24296 11936 24360 11940
rect 24376 11996 24440 12000
rect 24376 11940 24380 11996
rect 24380 11940 24436 11996
rect 24436 11940 24440 11996
rect 24376 11936 24440 11940
rect 24456 11996 24520 12000
rect 24456 11940 24460 11996
rect 24460 11940 24516 11996
rect 24516 11940 24520 11996
rect 24456 11936 24520 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 12216 11452 12280 11456
rect 12216 11396 12220 11452
rect 12220 11396 12276 11452
rect 12276 11396 12280 11452
rect 12216 11392 12280 11396
rect 12296 11452 12360 11456
rect 12296 11396 12300 11452
rect 12300 11396 12356 11452
rect 12356 11396 12360 11452
rect 12296 11392 12360 11396
rect 12376 11452 12440 11456
rect 12376 11396 12380 11452
rect 12380 11396 12436 11452
rect 12436 11396 12440 11452
rect 12376 11392 12440 11396
rect 12456 11452 12520 11456
rect 12456 11396 12460 11452
rect 12460 11396 12516 11452
rect 12516 11396 12520 11452
rect 12456 11392 12520 11396
rect 20216 11452 20280 11456
rect 20216 11396 20220 11452
rect 20220 11396 20276 11452
rect 20276 11396 20280 11452
rect 20216 11392 20280 11396
rect 20296 11452 20360 11456
rect 20296 11396 20300 11452
rect 20300 11396 20356 11452
rect 20356 11396 20360 11452
rect 20296 11392 20360 11396
rect 20376 11452 20440 11456
rect 20376 11396 20380 11452
rect 20380 11396 20436 11452
rect 20436 11396 20440 11452
rect 20376 11392 20440 11396
rect 20456 11452 20520 11456
rect 20456 11396 20460 11452
rect 20460 11396 20516 11452
rect 20516 11396 20520 11452
rect 20456 11392 20520 11396
rect 8216 10908 8280 10912
rect 8216 10852 8220 10908
rect 8220 10852 8276 10908
rect 8276 10852 8280 10908
rect 8216 10848 8280 10852
rect 8296 10908 8360 10912
rect 8296 10852 8300 10908
rect 8300 10852 8356 10908
rect 8356 10852 8360 10908
rect 8296 10848 8360 10852
rect 8376 10908 8440 10912
rect 8376 10852 8380 10908
rect 8380 10852 8436 10908
rect 8436 10852 8440 10908
rect 8376 10848 8440 10852
rect 8456 10908 8520 10912
rect 8456 10852 8460 10908
rect 8460 10852 8516 10908
rect 8516 10852 8520 10908
rect 8456 10848 8520 10852
rect 16216 10908 16280 10912
rect 16216 10852 16220 10908
rect 16220 10852 16276 10908
rect 16276 10852 16280 10908
rect 16216 10848 16280 10852
rect 16296 10908 16360 10912
rect 16296 10852 16300 10908
rect 16300 10852 16356 10908
rect 16356 10852 16360 10908
rect 16296 10848 16360 10852
rect 16376 10908 16440 10912
rect 16376 10852 16380 10908
rect 16380 10852 16436 10908
rect 16436 10852 16440 10908
rect 16376 10848 16440 10852
rect 16456 10908 16520 10912
rect 16456 10852 16460 10908
rect 16460 10852 16516 10908
rect 16516 10852 16520 10908
rect 16456 10848 16520 10852
rect 24216 10908 24280 10912
rect 24216 10852 24220 10908
rect 24220 10852 24276 10908
rect 24276 10852 24280 10908
rect 24216 10848 24280 10852
rect 24296 10908 24360 10912
rect 24296 10852 24300 10908
rect 24300 10852 24356 10908
rect 24356 10852 24360 10908
rect 24296 10848 24360 10852
rect 24376 10908 24440 10912
rect 24376 10852 24380 10908
rect 24380 10852 24436 10908
rect 24436 10852 24440 10908
rect 24376 10848 24440 10852
rect 24456 10908 24520 10912
rect 24456 10852 24460 10908
rect 24460 10852 24516 10908
rect 24516 10852 24520 10908
rect 24456 10848 24520 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 12216 10364 12280 10368
rect 12216 10308 12220 10364
rect 12220 10308 12276 10364
rect 12276 10308 12280 10364
rect 12216 10304 12280 10308
rect 12296 10364 12360 10368
rect 12296 10308 12300 10364
rect 12300 10308 12356 10364
rect 12356 10308 12360 10364
rect 12296 10304 12360 10308
rect 12376 10364 12440 10368
rect 12376 10308 12380 10364
rect 12380 10308 12436 10364
rect 12436 10308 12440 10364
rect 12376 10304 12440 10308
rect 12456 10364 12520 10368
rect 12456 10308 12460 10364
rect 12460 10308 12516 10364
rect 12516 10308 12520 10364
rect 12456 10304 12520 10308
rect 20216 10364 20280 10368
rect 20216 10308 20220 10364
rect 20220 10308 20276 10364
rect 20276 10308 20280 10364
rect 20216 10304 20280 10308
rect 20296 10364 20360 10368
rect 20296 10308 20300 10364
rect 20300 10308 20356 10364
rect 20356 10308 20360 10364
rect 20296 10304 20360 10308
rect 20376 10364 20440 10368
rect 20376 10308 20380 10364
rect 20380 10308 20436 10364
rect 20436 10308 20440 10364
rect 20376 10304 20440 10308
rect 20456 10364 20520 10368
rect 20456 10308 20460 10364
rect 20460 10308 20516 10364
rect 20516 10308 20520 10364
rect 20456 10304 20520 10308
rect 8216 9820 8280 9824
rect 8216 9764 8220 9820
rect 8220 9764 8276 9820
rect 8276 9764 8280 9820
rect 8216 9760 8280 9764
rect 8296 9820 8360 9824
rect 8296 9764 8300 9820
rect 8300 9764 8356 9820
rect 8356 9764 8360 9820
rect 8296 9760 8360 9764
rect 8376 9820 8440 9824
rect 8376 9764 8380 9820
rect 8380 9764 8436 9820
rect 8436 9764 8440 9820
rect 8376 9760 8440 9764
rect 8456 9820 8520 9824
rect 8456 9764 8460 9820
rect 8460 9764 8516 9820
rect 8516 9764 8520 9820
rect 8456 9760 8520 9764
rect 16216 9820 16280 9824
rect 16216 9764 16220 9820
rect 16220 9764 16276 9820
rect 16276 9764 16280 9820
rect 16216 9760 16280 9764
rect 16296 9820 16360 9824
rect 16296 9764 16300 9820
rect 16300 9764 16356 9820
rect 16356 9764 16360 9820
rect 16296 9760 16360 9764
rect 16376 9820 16440 9824
rect 16376 9764 16380 9820
rect 16380 9764 16436 9820
rect 16436 9764 16440 9820
rect 16376 9760 16440 9764
rect 16456 9820 16520 9824
rect 16456 9764 16460 9820
rect 16460 9764 16516 9820
rect 16516 9764 16520 9820
rect 16456 9760 16520 9764
rect 24216 9820 24280 9824
rect 24216 9764 24220 9820
rect 24220 9764 24276 9820
rect 24276 9764 24280 9820
rect 24216 9760 24280 9764
rect 24296 9820 24360 9824
rect 24296 9764 24300 9820
rect 24300 9764 24356 9820
rect 24356 9764 24360 9820
rect 24296 9760 24360 9764
rect 24376 9820 24440 9824
rect 24376 9764 24380 9820
rect 24380 9764 24436 9820
rect 24436 9764 24440 9820
rect 24376 9760 24440 9764
rect 24456 9820 24520 9824
rect 24456 9764 24460 9820
rect 24460 9764 24516 9820
rect 24516 9764 24520 9820
rect 24456 9760 24520 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 12216 9276 12280 9280
rect 12216 9220 12220 9276
rect 12220 9220 12276 9276
rect 12276 9220 12280 9276
rect 12216 9216 12280 9220
rect 12296 9276 12360 9280
rect 12296 9220 12300 9276
rect 12300 9220 12356 9276
rect 12356 9220 12360 9276
rect 12296 9216 12360 9220
rect 12376 9276 12440 9280
rect 12376 9220 12380 9276
rect 12380 9220 12436 9276
rect 12436 9220 12440 9276
rect 12376 9216 12440 9220
rect 12456 9276 12520 9280
rect 12456 9220 12460 9276
rect 12460 9220 12516 9276
rect 12516 9220 12520 9276
rect 12456 9216 12520 9220
rect 20216 9276 20280 9280
rect 20216 9220 20220 9276
rect 20220 9220 20276 9276
rect 20276 9220 20280 9276
rect 20216 9216 20280 9220
rect 20296 9276 20360 9280
rect 20296 9220 20300 9276
rect 20300 9220 20356 9276
rect 20356 9220 20360 9276
rect 20296 9216 20360 9220
rect 20376 9276 20440 9280
rect 20376 9220 20380 9276
rect 20380 9220 20436 9276
rect 20436 9220 20440 9276
rect 20376 9216 20440 9220
rect 20456 9276 20520 9280
rect 20456 9220 20460 9276
rect 20460 9220 20516 9276
rect 20516 9220 20520 9276
rect 20456 9216 20520 9220
rect 8216 8732 8280 8736
rect 8216 8676 8220 8732
rect 8220 8676 8276 8732
rect 8276 8676 8280 8732
rect 8216 8672 8280 8676
rect 8296 8732 8360 8736
rect 8296 8676 8300 8732
rect 8300 8676 8356 8732
rect 8356 8676 8360 8732
rect 8296 8672 8360 8676
rect 8376 8732 8440 8736
rect 8376 8676 8380 8732
rect 8380 8676 8436 8732
rect 8436 8676 8440 8732
rect 8376 8672 8440 8676
rect 8456 8732 8520 8736
rect 8456 8676 8460 8732
rect 8460 8676 8516 8732
rect 8516 8676 8520 8732
rect 8456 8672 8520 8676
rect 16216 8732 16280 8736
rect 16216 8676 16220 8732
rect 16220 8676 16276 8732
rect 16276 8676 16280 8732
rect 16216 8672 16280 8676
rect 16296 8732 16360 8736
rect 16296 8676 16300 8732
rect 16300 8676 16356 8732
rect 16356 8676 16360 8732
rect 16296 8672 16360 8676
rect 16376 8732 16440 8736
rect 16376 8676 16380 8732
rect 16380 8676 16436 8732
rect 16436 8676 16440 8732
rect 16376 8672 16440 8676
rect 16456 8732 16520 8736
rect 16456 8676 16460 8732
rect 16460 8676 16516 8732
rect 16516 8676 16520 8732
rect 16456 8672 16520 8676
rect 24216 8732 24280 8736
rect 24216 8676 24220 8732
rect 24220 8676 24276 8732
rect 24276 8676 24280 8732
rect 24216 8672 24280 8676
rect 24296 8732 24360 8736
rect 24296 8676 24300 8732
rect 24300 8676 24356 8732
rect 24356 8676 24360 8732
rect 24296 8672 24360 8676
rect 24376 8732 24440 8736
rect 24376 8676 24380 8732
rect 24380 8676 24436 8732
rect 24436 8676 24440 8732
rect 24376 8672 24440 8676
rect 24456 8732 24520 8736
rect 24456 8676 24460 8732
rect 24460 8676 24516 8732
rect 24516 8676 24520 8732
rect 24456 8672 24520 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 12216 8188 12280 8192
rect 12216 8132 12220 8188
rect 12220 8132 12276 8188
rect 12276 8132 12280 8188
rect 12216 8128 12280 8132
rect 12296 8188 12360 8192
rect 12296 8132 12300 8188
rect 12300 8132 12356 8188
rect 12356 8132 12360 8188
rect 12296 8128 12360 8132
rect 12376 8188 12440 8192
rect 12376 8132 12380 8188
rect 12380 8132 12436 8188
rect 12436 8132 12440 8188
rect 12376 8128 12440 8132
rect 12456 8188 12520 8192
rect 12456 8132 12460 8188
rect 12460 8132 12516 8188
rect 12516 8132 12520 8188
rect 12456 8128 12520 8132
rect 20216 8188 20280 8192
rect 20216 8132 20220 8188
rect 20220 8132 20276 8188
rect 20276 8132 20280 8188
rect 20216 8128 20280 8132
rect 20296 8188 20360 8192
rect 20296 8132 20300 8188
rect 20300 8132 20356 8188
rect 20356 8132 20360 8188
rect 20296 8128 20360 8132
rect 20376 8188 20440 8192
rect 20376 8132 20380 8188
rect 20380 8132 20436 8188
rect 20436 8132 20440 8188
rect 20376 8128 20440 8132
rect 20456 8188 20520 8192
rect 20456 8132 20460 8188
rect 20460 8132 20516 8188
rect 20516 8132 20520 8188
rect 20456 8128 20520 8132
rect 8216 7644 8280 7648
rect 8216 7588 8220 7644
rect 8220 7588 8276 7644
rect 8276 7588 8280 7644
rect 8216 7584 8280 7588
rect 8296 7644 8360 7648
rect 8296 7588 8300 7644
rect 8300 7588 8356 7644
rect 8356 7588 8360 7644
rect 8296 7584 8360 7588
rect 8376 7644 8440 7648
rect 8376 7588 8380 7644
rect 8380 7588 8436 7644
rect 8436 7588 8440 7644
rect 8376 7584 8440 7588
rect 8456 7644 8520 7648
rect 8456 7588 8460 7644
rect 8460 7588 8516 7644
rect 8516 7588 8520 7644
rect 8456 7584 8520 7588
rect 16216 7644 16280 7648
rect 16216 7588 16220 7644
rect 16220 7588 16276 7644
rect 16276 7588 16280 7644
rect 16216 7584 16280 7588
rect 16296 7644 16360 7648
rect 16296 7588 16300 7644
rect 16300 7588 16356 7644
rect 16356 7588 16360 7644
rect 16296 7584 16360 7588
rect 16376 7644 16440 7648
rect 16376 7588 16380 7644
rect 16380 7588 16436 7644
rect 16436 7588 16440 7644
rect 16376 7584 16440 7588
rect 16456 7644 16520 7648
rect 16456 7588 16460 7644
rect 16460 7588 16516 7644
rect 16516 7588 16520 7644
rect 16456 7584 16520 7588
rect 24216 7644 24280 7648
rect 24216 7588 24220 7644
rect 24220 7588 24276 7644
rect 24276 7588 24280 7644
rect 24216 7584 24280 7588
rect 24296 7644 24360 7648
rect 24296 7588 24300 7644
rect 24300 7588 24356 7644
rect 24356 7588 24360 7644
rect 24296 7584 24360 7588
rect 24376 7644 24440 7648
rect 24376 7588 24380 7644
rect 24380 7588 24436 7644
rect 24436 7588 24440 7644
rect 24376 7584 24440 7588
rect 24456 7644 24520 7648
rect 24456 7588 24460 7644
rect 24460 7588 24516 7644
rect 24516 7588 24520 7644
rect 24456 7584 24520 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 12216 7100 12280 7104
rect 12216 7044 12220 7100
rect 12220 7044 12276 7100
rect 12276 7044 12280 7100
rect 12216 7040 12280 7044
rect 12296 7100 12360 7104
rect 12296 7044 12300 7100
rect 12300 7044 12356 7100
rect 12356 7044 12360 7100
rect 12296 7040 12360 7044
rect 12376 7100 12440 7104
rect 12376 7044 12380 7100
rect 12380 7044 12436 7100
rect 12436 7044 12440 7100
rect 12376 7040 12440 7044
rect 12456 7100 12520 7104
rect 12456 7044 12460 7100
rect 12460 7044 12516 7100
rect 12516 7044 12520 7100
rect 12456 7040 12520 7044
rect 20216 7100 20280 7104
rect 20216 7044 20220 7100
rect 20220 7044 20276 7100
rect 20276 7044 20280 7100
rect 20216 7040 20280 7044
rect 20296 7100 20360 7104
rect 20296 7044 20300 7100
rect 20300 7044 20356 7100
rect 20356 7044 20360 7100
rect 20296 7040 20360 7044
rect 20376 7100 20440 7104
rect 20376 7044 20380 7100
rect 20380 7044 20436 7100
rect 20436 7044 20440 7100
rect 20376 7040 20440 7044
rect 20456 7100 20520 7104
rect 20456 7044 20460 7100
rect 20460 7044 20516 7100
rect 20516 7044 20520 7100
rect 20456 7040 20520 7044
rect 8216 6556 8280 6560
rect 8216 6500 8220 6556
rect 8220 6500 8276 6556
rect 8276 6500 8280 6556
rect 8216 6496 8280 6500
rect 8296 6556 8360 6560
rect 8296 6500 8300 6556
rect 8300 6500 8356 6556
rect 8356 6500 8360 6556
rect 8296 6496 8360 6500
rect 8376 6556 8440 6560
rect 8376 6500 8380 6556
rect 8380 6500 8436 6556
rect 8436 6500 8440 6556
rect 8376 6496 8440 6500
rect 8456 6556 8520 6560
rect 8456 6500 8460 6556
rect 8460 6500 8516 6556
rect 8516 6500 8520 6556
rect 8456 6496 8520 6500
rect 16216 6556 16280 6560
rect 16216 6500 16220 6556
rect 16220 6500 16276 6556
rect 16276 6500 16280 6556
rect 16216 6496 16280 6500
rect 16296 6556 16360 6560
rect 16296 6500 16300 6556
rect 16300 6500 16356 6556
rect 16356 6500 16360 6556
rect 16296 6496 16360 6500
rect 16376 6556 16440 6560
rect 16376 6500 16380 6556
rect 16380 6500 16436 6556
rect 16436 6500 16440 6556
rect 16376 6496 16440 6500
rect 16456 6556 16520 6560
rect 16456 6500 16460 6556
rect 16460 6500 16516 6556
rect 16516 6500 16520 6556
rect 16456 6496 16520 6500
rect 24216 6556 24280 6560
rect 24216 6500 24220 6556
rect 24220 6500 24276 6556
rect 24276 6500 24280 6556
rect 24216 6496 24280 6500
rect 24296 6556 24360 6560
rect 24296 6500 24300 6556
rect 24300 6500 24356 6556
rect 24356 6500 24360 6556
rect 24296 6496 24360 6500
rect 24376 6556 24440 6560
rect 24376 6500 24380 6556
rect 24380 6500 24436 6556
rect 24436 6500 24440 6556
rect 24376 6496 24440 6500
rect 24456 6556 24520 6560
rect 24456 6500 24460 6556
rect 24460 6500 24516 6556
rect 24516 6500 24520 6556
rect 24456 6496 24520 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 12216 6012 12280 6016
rect 12216 5956 12220 6012
rect 12220 5956 12276 6012
rect 12276 5956 12280 6012
rect 12216 5952 12280 5956
rect 12296 6012 12360 6016
rect 12296 5956 12300 6012
rect 12300 5956 12356 6012
rect 12356 5956 12360 6012
rect 12296 5952 12360 5956
rect 12376 6012 12440 6016
rect 12376 5956 12380 6012
rect 12380 5956 12436 6012
rect 12436 5956 12440 6012
rect 12376 5952 12440 5956
rect 12456 6012 12520 6016
rect 12456 5956 12460 6012
rect 12460 5956 12516 6012
rect 12516 5956 12520 6012
rect 12456 5952 12520 5956
rect 20216 6012 20280 6016
rect 20216 5956 20220 6012
rect 20220 5956 20276 6012
rect 20276 5956 20280 6012
rect 20216 5952 20280 5956
rect 20296 6012 20360 6016
rect 20296 5956 20300 6012
rect 20300 5956 20356 6012
rect 20356 5956 20360 6012
rect 20296 5952 20360 5956
rect 20376 6012 20440 6016
rect 20376 5956 20380 6012
rect 20380 5956 20436 6012
rect 20436 5956 20440 6012
rect 20376 5952 20440 5956
rect 20456 6012 20520 6016
rect 20456 5956 20460 6012
rect 20460 5956 20516 6012
rect 20516 5956 20520 6012
rect 20456 5952 20520 5956
rect 8216 5468 8280 5472
rect 8216 5412 8220 5468
rect 8220 5412 8276 5468
rect 8276 5412 8280 5468
rect 8216 5408 8280 5412
rect 8296 5468 8360 5472
rect 8296 5412 8300 5468
rect 8300 5412 8356 5468
rect 8356 5412 8360 5468
rect 8296 5408 8360 5412
rect 8376 5468 8440 5472
rect 8376 5412 8380 5468
rect 8380 5412 8436 5468
rect 8436 5412 8440 5468
rect 8376 5408 8440 5412
rect 8456 5468 8520 5472
rect 8456 5412 8460 5468
rect 8460 5412 8516 5468
rect 8516 5412 8520 5468
rect 8456 5408 8520 5412
rect 16216 5468 16280 5472
rect 16216 5412 16220 5468
rect 16220 5412 16276 5468
rect 16276 5412 16280 5468
rect 16216 5408 16280 5412
rect 16296 5468 16360 5472
rect 16296 5412 16300 5468
rect 16300 5412 16356 5468
rect 16356 5412 16360 5468
rect 16296 5408 16360 5412
rect 16376 5468 16440 5472
rect 16376 5412 16380 5468
rect 16380 5412 16436 5468
rect 16436 5412 16440 5468
rect 16376 5408 16440 5412
rect 16456 5468 16520 5472
rect 16456 5412 16460 5468
rect 16460 5412 16516 5468
rect 16516 5412 16520 5468
rect 16456 5408 16520 5412
rect 24216 5468 24280 5472
rect 24216 5412 24220 5468
rect 24220 5412 24276 5468
rect 24276 5412 24280 5468
rect 24216 5408 24280 5412
rect 24296 5468 24360 5472
rect 24296 5412 24300 5468
rect 24300 5412 24356 5468
rect 24356 5412 24360 5468
rect 24296 5408 24360 5412
rect 24376 5468 24440 5472
rect 24376 5412 24380 5468
rect 24380 5412 24436 5468
rect 24436 5412 24440 5468
rect 24376 5408 24440 5412
rect 24456 5468 24520 5472
rect 24456 5412 24460 5468
rect 24460 5412 24516 5468
rect 24516 5412 24520 5468
rect 24456 5408 24520 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 12216 4924 12280 4928
rect 12216 4868 12220 4924
rect 12220 4868 12276 4924
rect 12276 4868 12280 4924
rect 12216 4864 12280 4868
rect 12296 4924 12360 4928
rect 12296 4868 12300 4924
rect 12300 4868 12356 4924
rect 12356 4868 12360 4924
rect 12296 4864 12360 4868
rect 12376 4924 12440 4928
rect 12376 4868 12380 4924
rect 12380 4868 12436 4924
rect 12436 4868 12440 4924
rect 12376 4864 12440 4868
rect 12456 4924 12520 4928
rect 12456 4868 12460 4924
rect 12460 4868 12516 4924
rect 12516 4868 12520 4924
rect 12456 4864 12520 4868
rect 20216 4924 20280 4928
rect 20216 4868 20220 4924
rect 20220 4868 20276 4924
rect 20276 4868 20280 4924
rect 20216 4864 20280 4868
rect 20296 4924 20360 4928
rect 20296 4868 20300 4924
rect 20300 4868 20356 4924
rect 20356 4868 20360 4924
rect 20296 4864 20360 4868
rect 20376 4924 20440 4928
rect 20376 4868 20380 4924
rect 20380 4868 20436 4924
rect 20436 4868 20440 4924
rect 20376 4864 20440 4868
rect 20456 4924 20520 4928
rect 20456 4868 20460 4924
rect 20460 4868 20516 4924
rect 20516 4868 20520 4924
rect 20456 4864 20520 4868
rect 8216 4380 8280 4384
rect 8216 4324 8220 4380
rect 8220 4324 8276 4380
rect 8276 4324 8280 4380
rect 8216 4320 8280 4324
rect 8296 4380 8360 4384
rect 8296 4324 8300 4380
rect 8300 4324 8356 4380
rect 8356 4324 8360 4380
rect 8296 4320 8360 4324
rect 8376 4380 8440 4384
rect 8376 4324 8380 4380
rect 8380 4324 8436 4380
rect 8436 4324 8440 4380
rect 8376 4320 8440 4324
rect 8456 4380 8520 4384
rect 8456 4324 8460 4380
rect 8460 4324 8516 4380
rect 8516 4324 8520 4380
rect 8456 4320 8520 4324
rect 16216 4380 16280 4384
rect 16216 4324 16220 4380
rect 16220 4324 16276 4380
rect 16276 4324 16280 4380
rect 16216 4320 16280 4324
rect 16296 4380 16360 4384
rect 16296 4324 16300 4380
rect 16300 4324 16356 4380
rect 16356 4324 16360 4380
rect 16296 4320 16360 4324
rect 16376 4380 16440 4384
rect 16376 4324 16380 4380
rect 16380 4324 16436 4380
rect 16436 4324 16440 4380
rect 16376 4320 16440 4324
rect 16456 4380 16520 4384
rect 16456 4324 16460 4380
rect 16460 4324 16516 4380
rect 16516 4324 16520 4380
rect 16456 4320 16520 4324
rect 24216 4380 24280 4384
rect 24216 4324 24220 4380
rect 24220 4324 24276 4380
rect 24276 4324 24280 4380
rect 24216 4320 24280 4324
rect 24296 4380 24360 4384
rect 24296 4324 24300 4380
rect 24300 4324 24356 4380
rect 24356 4324 24360 4380
rect 24296 4320 24360 4324
rect 24376 4380 24440 4384
rect 24376 4324 24380 4380
rect 24380 4324 24436 4380
rect 24436 4324 24440 4380
rect 24376 4320 24440 4324
rect 24456 4380 24520 4384
rect 24456 4324 24460 4380
rect 24460 4324 24516 4380
rect 24516 4324 24520 4380
rect 24456 4320 24520 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 12216 3836 12280 3840
rect 12216 3780 12220 3836
rect 12220 3780 12276 3836
rect 12276 3780 12280 3836
rect 12216 3776 12280 3780
rect 12296 3836 12360 3840
rect 12296 3780 12300 3836
rect 12300 3780 12356 3836
rect 12356 3780 12360 3836
rect 12296 3776 12360 3780
rect 12376 3836 12440 3840
rect 12376 3780 12380 3836
rect 12380 3780 12436 3836
rect 12436 3780 12440 3836
rect 12376 3776 12440 3780
rect 12456 3836 12520 3840
rect 12456 3780 12460 3836
rect 12460 3780 12516 3836
rect 12516 3780 12520 3836
rect 12456 3776 12520 3780
rect 20216 3836 20280 3840
rect 20216 3780 20220 3836
rect 20220 3780 20276 3836
rect 20276 3780 20280 3836
rect 20216 3776 20280 3780
rect 20296 3836 20360 3840
rect 20296 3780 20300 3836
rect 20300 3780 20356 3836
rect 20356 3780 20360 3836
rect 20296 3776 20360 3780
rect 20376 3836 20440 3840
rect 20376 3780 20380 3836
rect 20380 3780 20436 3836
rect 20436 3780 20440 3836
rect 20376 3776 20440 3780
rect 20456 3836 20520 3840
rect 20456 3780 20460 3836
rect 20460 3780 20516 3836
rect 20516 3780 20520 3836
rect 20456 3776 20520 3780
rect 8216 3292 8280 3296
rect 8216 3236 8220 3292
rect 8220 3236 8276 3292
rect 8276 3236 8280 3292
rect 8216 3232 8280 3236
rect 8296 3292 8360 3296
rect 8296 3236 8300 3292
rect 8300 3236 8356 3292
rect 8356 3236 8360 3292
rect 8296 3232 8360 3236
rect 8376 3292 8440 3296
rect 8376 3236 8380 3292
rect 8380 3236 8436 3292
rect 8436 3236 8440 3292
rect 8376 3232 8440 3236
rect 8456 3292 8520 3296
rect 8456 3236 8460 3292
rect 8460 3236 8516 3292
rect 8516 3236 8520 3292
rect 8456 3232 8520 3236
rect 16216 3292 16280 3296
rect 16216 3236 16220 3292
rect 16220 3236 16276 3292
rect 16276 3236 16280 3292
rect 16216 3232 16280 3236
rect 16296 3292 16360 3296
rect 16296 3236 16300 3292
rect 16300 3236 16356 3292
rect 16356 3236 16360 3292
rect 16296 3232 16360 3236
rect 16376 3292 16440 3296
rect 16376 3236 16380 3292
rect 16380 3236 16436 3292
rect 16436 3236 16440 3292
rect 16376 3232 16440 3236
rect 16456 3292 16520 3296
rect 16456 3236 16460 3292
rect 16460 3236 16516 3292
rect 16516 3236 16520 3292
rect 16456 3232 16520 3236
rect 24216 3292 24280 3296
rect 24216 3236 24220 3292
rect 24220 3236 24276 3292
rect 24276 3236 24280 3292
rect 24216 3232 24280 3236
rect 24296 3292 24360 3296
rect 24296 3236 24300 3292
rect 24300 3236 24356 3292
rect 24356 3236 24360 3292
rect 24296 3232 24360 3236
rect 24376 3292 24440 3296
rect 24376 3236 24380 3292
rect 24380 3236 24436 3292
rect 24436 3236 24440 3292
rect 24376 3232 24440 3236
rect 24456 3292 24520 3296
rect 24456 3236 24460 3292
rect 24460 3236 24516 3292
rect 24516 3236 24520 3292
rect 24456 3232 24520 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 12216 2748 12280 2752
rect 12216 2692 12220 2748
rect 12220 2692 12276 2748
rect 12276 2692 12280 2748
rect 12216 2688 12280 2692
rect 12296 2748 12360 2752
rect 12296 2692 12300 2748
rect 12300 2692 12356 2748
rect 12356 2692 12360 2748
rect 12296 2688 12360 2692
rect 12376 2748 12440 2752
rect 12376 2692 12380 2748
rect 12380 2692 12436 2748
rect 12436 2692 12440 2748
rect 12376 2688 12440 2692
rect 12456 2748 12520 2752
rect 12456 2692 12460 2748
rect 12460 2692 12516 2748
rect 12516 2692 12520 2748
rect 12456 2688 12520 2692
rect 20216 2748 20280 2752
rect 20216 2692 20220 2748
rect 20220 2692 20276 2748
rect 20276 2692 20280 2748
rect 20216 2688 20280 2692
rect 20296 2748 20360 2752
rect 20296 2692 20300 2748
rect 20300 2692 20356 2748
rect 20356 2692 20360 2748
rect 20296 2688 20360 2692
rect 20376 2748 20440 2752
rect 20376 2692 20380 2748
rect 20380 2692 20436 2748
rect 20436 2692 20440 2748
rect 20376 2688 20440 2692
rect 20456 2748 20520 2752
rect 20456 2692 20460 2748
rect 20460 2692 20516 2748
rect 20516 2692 20520 2748
rect 20456 2688 20520 2692
rect 8216 2204 8280 2208
rect 8216 2148 8220 2204
rect 8220 2148 8276 2204
rect 8276 2148 8280 2204
rect 8216 2144 8280 2148
rect 8296 2204 8360 2208
rect 8296 2148 8300 2204
rect 8300 2148 8356 2204
rect 8356 2148 8360 2204
rect 8296 2144 8360 2148
rect 8376 2204 8440 2208
rect 8376 2148 8380 2204
rect 8380 2148 8436 2204
rect 8436 2148 8440 2204
rect 8376 2144 8440 2148
rect 8456 2204 8520 2208
rect 8456 2148 8460 2204
rect 8460 2148 8516 2204
rect 8516 2148 8520 2204
rect 8456 2144 8520 2148
rect 16216 2204 16280 2208
rect 16216 2148 16220 2204
rect 16220 2148 16276 2204
rect 16276 2148 16280 2204
rect 16216 2144 16280 2148
rect 16296 2204 16360 2208
rect 16296 2148 16300 2204
rect 16300 2148 16356 2204
rect 16356 2148 16360 2204
rect 16296 2144 16360 2148
rect 16376 2204 16440 2208
rect 16376 2148 16380 2204
rect 16380 2148 16436 2204
rect 16436 2148 16440 2204
rect 16376 2144 16440 2148
rect 16456 2204 16520 2208
rect 16456 2148 16460 2204
rect 16460 2148 16516 2204
rect 16516 2148 16520 2204
rect 16456 2144 16520 2148
rect 24216 2204 24280 2208
rect 24216 2148 24220 2204
rect 24220 2148 24276 2204
rect 24276 2148 24280 2204
rect 24216 2144 24280 2148
rect 24296 2204 24360 2208
rect 24296 2148 24300 2204
rect 24300 2148 24356 2204
rect 24356 2148 24360 2204
rect 24296 2144 24360 2148
rect 24376 2204 24440 2208
rect 24376 2148 24380 2204
rect 24380 2148 24436 2204
rect 24436 2148 24440 2204
rect 24376 2144 24440 2148
rect 24456 2204 24520 2208
rect 24456 2148 24460 2204
rect 24460 2148 24516 2204
rect 24516 2148 24520 2204
rect 24456 2144 24520 2148
rect 4216 1660 4280 1664
rect 4216 1604 4220 1660
rect 4220 1604 4276 1660
rect 4276 1604 4280 1660
rect 4216 1600 4280 1604
rect 4296 1660 4360 1664
rect 4296 1604 4300 1660
rect 4300 1604 4356 1660
rect 4356 1604 4360 1660
rect 4296 1600 4360 1604
rect 4376 1660 4440 1664
rect 4376 1604 4380 1660
rect 4380 1604 4436 1660
rect 4436 1604 4440 1660
rect 4376 1600 4440 1604
rect 4456 1660 4520 1664
rect 4456 1604 4460 1660
rect 4460 1604 4516 1660
rect 4516 1604 4520 1660
rect 4456 1600 4520 1604
rect 12216 1660 12280 1664
rect 12216 1604 12220 1660
rect 12220 1604 12276 1660
rect 12276 1604 12280 1660
rect 12216 1600 12280 1604
rect 12296 1660 12360 1664
rect 12296 1604 12300 1660
rect 12300 1604 12356 1660
rect 12356 1604 12360 1660
rect 12296 1600 12360 1604
rect 12376 1660 12440 1664
rect 12376 1604 12380 1660
rect 12380 1604 12436 1660
rect 12436 1604 12440 1660
rect 12376 1600 12440 1604
rect 12456 1660 12520 1664
rect 12456 1604 12460 1660
rect 12460 1604 12516 1660
rect 12516 1604 12520 1660
rect 12456 1600 12520 1604
rect 20216 1660 20280 1664
rect 20216 1604 20220 1660
rect 20220 1604 20276 1660
rect 20276 1604 20280 1660
rect 20216 1600 20280 1604
rect 20296 1660 20360 1664
rect 20296 1604 20300 1660
rect 20300 1604 20356 1660
rect 20356 1604 20360 1660
rect 20296 1600 20360 1604
rect 20376 1660 20440 1664
rect 20376 1604 20380 1660
rect 20380 1604 20436 1660
rect 20436 1604 20440 1660
rect 20376 1600 20440 1604
rect 20456 1660 20520 1664
rect 20456 1604 20460 1660
rect 20460 1604 20516 1660
rect 20516 1604 20520 1660
rect 20456 1600 20520 1604
rect 8216 1116 8280 1120
rect 8216 1060 8220 1116
rect 8220 1060 8276 1116
rect 8276 1060 8280 1116
rect 8216 1056 8280 1060
rect 8296 1116 8360 1120
rect 8296 1060 8300 1116
rect 8300 1060 8356 1116
rect 8356 1060 8360 1116
rect 8296 1056 8360 1060
rect 8376 1116 8440 1120
rect 8376 1060 8380 1116
rect 8380 1060 8436 1116
rect 8436 1060 8440 1116
rect 8376 1056 8440 1060
rect 8456 1116 8520 1120
rect 8456 1060 8460 1116
rect 8460 1060 8516 1116
rect 8516 1060 8520 1116
rect 8456 1056 8520 1060
rect 16216 1116 16280 1120
rect 16216 1060 16220 1116
rect 16220 1060 16276 1116
rect 16276 1060 16280 1116
rect 16216 1056 16280 1060
rect 16296 1116 16360 1120
rect 16296 1060 16300 1116
rect 16300 1060 16356 1116
rect 16356 1060 16360 1116
rect 16296 1056 16360 1060
rect 16376 1116 16440 1120
rect 16376 1060 16380 1116
rect 16380 1060 16436 1116
rect 16436 1060 16440 1116
rect 16376 1056 16440 1060
rect 16456 1116 16520 1120
rect 16456 1060 16460 1116
rect 16460 1060 16516 1116
rect 16516 1060 16520 1116
rect 16456 1056 16520 1060
rect 24216 1116 24280 1120
rect 24216 1060 24220 1116
rect 24220 1060 24276 1116
rect 24276 1060 24280 1116
rect 24216 1056 24280 1060
rect 24296 1116 24360 1120
rect 24296 1060 24300 1116
rect 24300 1060 24356 1116
rect 24356 1060 24360 1116
rect 24296 1056 24360 1060
rect 24376 1116 24440 1120
rect 24376 1060 24380 1116
rect 24380 1060 24436 1116
rect 24436 1060 24440 1116
rect 24376 1056 24440 1060
rect 24456 1116 24520 1120
rect 24456 1060 24460 1116
rect 24460 1060 24516 1116
rect 24516 1060 24520 1116
rect 24456 1056 24520 1060
<< metal4 >>
rect 4208 20160 4528 20720
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 1664 4528 2688
rect 4208 1600 4216 1664
rect 4280 1600 4296 1664
rect 4360 1600 4376 1664
rect 4440 1600 4456 1664
rect 4520 1600 4528 1664
rect 4208 1040 4528 1600
rect 8208 20704 8528 20720
rect 8208 20640 8216 20704
rect 8280 20640 8296 20704
rect 8360 20640 8376 20704
rect 8440 20640 8456 20704
rect 8520 20640 8528 20704
rect 8208 19616 8528 20640
rect 8208 19552 8216 19616
rect 8280 19552 8296 19616
rect 8360 19552 8376 19616
rect 8440 19552 8456 19616
rect 8520 19552 8528 19616
rect 8208 18528 8528 19552
rect 12208 20160 12528 20720
rect 12208 20096 12216 20160
rect 12280 20096 12296 20160
rect 12360 20096 12376 20160
rect 12440 20096 12456 20160
rect 12520 20096 12528 20160
rect 11467 19140 11533 19141
rect 11467 19076 11468 19140
rect 11532 19076 11533 19140
rect 11467 19075 11533 19076
rect 8208 18464 8216 18528
rect 8280 18464 8296 18528
rect 8360 18464 8376 18528
rect 8440 18464 8456 18528
rect 8520 18464 8528 18528
rect 8208 17440 8528 18464
rect 11470 17917 11530 19075
rect 12208 19072 12528 20096
rect 12208 19008 12216 19072
rect 12280 19008 12296 19072
rect 12360 19008 12376 19072
rect 12440 19008 12456 19072
rect 12520 19008 12528 19072
rect 11651 18868 11717 18869
rect 11651 18804 11652 18868
rect 11716 18804 11717 18868
rect 11651 18803 11717 18804
rect 11467 17916 11533 17917
rect 11467 17852 11468 17916
rect 11532 17852 11533 17916
rect 11467 17851 11533 17852
rect 8208 17376 8216 17440
rect 8280 17376 8296 17440
rect 8360 17376 8376 17440
rect 8440 17376 8456 17440
rect 8520 17376 8528 17440
rect 8208 16352 8528 17376
rect 8208 16288 8216 16352
rect 8280 16288 8296 16352
rect 8360 16288 8376 16352
rect 8440 16288 8456 16352
rect 8520 16288 8528 16352
rect 8208 15264 8528 16288
rect 11654 16285 11714 18803
rect 12208 17984 12528 19008
rect 12208 17920 12216 17984
rect 12280 17920 12296 17984
rect 12360 17920 12376 17984
rect 12440 17920 12456 17984
rect 12520 17920 12528 17984
rect 12208 16896 12528 17920
rect 12208 16832 12216 16896
rect 12280 16832 12296 16896
rect 12360 16832 12376 16896
rect 12440 16832 12456 16896
rect 12520 16832 12528 16896
rect 11651 16284 11717 16285
rect 11651 16220 11652 16284
rect 11716 16220 11717 16284
rect 11651 16219 11717 16220
rect 8208 15200 8216 15264
rect 8280 15200 8296 15264
rect 8360 15200 8376 15264
rect 8440 15200 8456 15264
rect 8520 15200 8528 15264
rect 8208 14176 8528 15200
rect 8208 14112 8216 14176
rect 8280 14112 8296 14176
rect 8360 14112 8376 14176
rect 8440 14112 8456 14176
rect 8520 14112 8528 14176
rect 8208 13088 8528 14112
rect 8208 13024 8216 13088
rect 8280 13024 8296 13088
rect 8360 13024 8376 13088
rect 8440 13024 8456 13088
rect 8520 13024 8528 13088
rect 8208 12000 8528 13024
rect 8208 11936 8216 12000
rect 8280 11936 8296 12000
rect 8360 11936 8376 12000
rect 8440 11936 8456 12000
rect 8520 11936 8528 12000
rect 8208 10912 8528 11936
rect 8208 10848 8216 10912
rect 8280 10848 8296 10912
rect 8360 10848 8376 10912
rect 8440 10848 8456 10912
rect 8520 10848 8528 10912
rect 8208 9824 8528 10848
rect 8208 9760 8216 9824
rect 8280 9760 8296 9824
rect 8360 9760 8376 9824
rect 8440 9760 8456 9824
rect 8520 9760 8528 9824
rect 8208 8736 8528 9760
rect 8208 8672 8216 8736
rect 8280 8672 8296 8736
rect 8360 8672 8376 8736
rect 8440 8672 8456 8736
rect 8520 8672 8528 8736
rect 8208 7648 8528 8672
rect 8208 7584 8216 7648
rect 8280 7584 8296 7648
rect 8360 7584 8376 7648
rect 8440 7584 8456 7648
rect 8520 7584 8528 7648
rect 8208 6560 8528 7584
rect 8208 6496 8216 6560
rect 8280 6496 8296 6560
rect 8360 6496 8376 6560
rect 8440 6496 8456 6560
rect 8520 6496 8528 6560
rect 8208 5472 8528 6496
rect 8208 5408 8216 5472
rect 8280 5408 8296 5472
rect 8360 5408 8376 5472
rect 8440 5408 8456 5472
rect 8520 5408 8528 5472
rect 8208 4384 8528 5408
rect 8208 4320 8216 4384
rect 8280 4320 8296 4384
rect 8360 4320 8376 4384
rect 8440 4320 8456 4384
rect 8520 4320 8528 4384
rect 8208 3296 8528 4320
rect 8208 3232 8216 3296
rect 8280 3232 8296 3296
rect 8360 3232 8376 3296
rect 8440 3232 8456 3296
rect 8520 3232 8528 3296
rect 8208 2208 8528 3232
rect 8208 2144 8216 2208
rect 8280 2144 8296 2208
rect 8360 2144 8376 2208
rect 8440 2144 8456 2208
rect 8520 2144 8528 2208
rect 8208 1120 8528 2144
rect 8208 1056 8216 1120
rect 8280 1056 8296 1120
rect 8360 1056 8376 1120
rect 8440 1056 8456 1120
rect 8520 1056 8528 1120
rect 8208 1040 8528 1056
rect 12208 15808 12528 16832
rect 12208 15744 12216 15808
rect 12280 15744 12296 15808
rect 12360 15744 12376 15808
rect 12440 15744 12456 15808
rect 12520 15744 12528 15808
rect 12208 14720 12528 15744
rect 12208 14656 12216 14720
rect 12280 14656 12296 14720
rect 12360 14656 12376 14720
rect 12440 14656 12456 14720
rect 12520 14656 12528 14720
rect 12208 13632 12528 14656
rect 12208 13568 12216 13632
rect 12280 13568 12296 13632
rect 12360 13568 12376 13632
rect 12440 13568 12456 13632
rect 12520 13568 12528 13632
rect 12208 12544 12528 13568
rect 12208 12480 12216 12544
rect 12280 12480 12296 12544
rect 12360 12480 12376 12544
rect 12440 12480 12456 12544
rect 12520 12480 12528 12544
rect 12208 11456 12528 12480
rect 12208 11392 12216 11456
rect 12280 11392 12296 11456
rect 12360 11392 12376 11456
rect 12440 11392 12456 11456
rect 12520 11392 12528 11456
rect 12208 10368 12528 11392
rect 12208 10304 12216 10368
rect 12280 10304 12296 10368
rect 12360 10304 12376 10368
rect 12440 10304 12456 10368
rect 12520 10304 12528 10368
rect 12208 9280 12528 10304
rect 12208 9216 12216 9280
rect 12280 9216 12296 9280
rect 12360 9216 12376 9280
rect 12440 9216 12456 9280
rect 12520 9216 12528 9280
rect 12208 8192 12528 9216
rect 12208 8128 12216 8192
rect 12280 8128 12296 8192
rect 12360 8128 12376 8192
rect 12440 8128 12456 8192
rect 12520 8128 12528 8192
rect 12208 7104 12528 8128
rect 12208 7040 12216 7104
rect 12280 7040 12296 7104
rect 12360 7040 12376 7104
rect 12440 7040 12456 7104
rect 12520 7040 12528 7104
rect 12208 6016 12528 7040
rect 12208 5952 12216 6016
rect 12280 5952 12296 6016
rect 12360 5952 12376 6016
rect 12440 5952 12456 6016
rect 12520 5952 12528 6016
rect 12208 4928 12528 5952
rect 12208 4864 12216 4928
rect 12280 4864 12296 4928
rect 12360 4864 12376 4928
rect 12440 4864 12456 4928
rect 12520 4864 12528 4928
rect 12208 3840 12528 4864
rect 12208 3776 12216 3840
rect 12280 3776 12296 3840
rect 12360 3776 12376 3840
rect 12440 3776 12456 3840
rect 12520 3776 12528 3840
rect 12208 2752 12528 3776
rect 12208 2688 12216 2752
rect 12280 2688 12296 2752
rect 12360 2688 12376 2752
rect 12440 2688 12456 2752
rect 12520 2688 12528 2752
rect 12208 1664 12528 2688
rect 12208 1600 12216 1664
rect 12280 1600 12296 1664
rect 12360 1600 12376 1664
rect 12440 1600 12456 1664
rect 12520 1600 12528 1664
rect 12208 1040 12528 1600
rect 16208 20704 16528 20720
rect 16208 20640 16216 20704
rect 16280 20640 16296 20704
rect 16360 20640 16376 20704
rect 16440 20640 16456 20704
rect 16520 20640 16528 20704
rect 16208 19616 16528 20640
rect 16208 19552 16216 19616
rect 16280 19552 16296 19616
rect 16360 19552 16376 19616
rect 16440 19552 16456 19616
rect 16520 19552 16528 19616
rect 16208 18528 16528 19552
rect 16208 18464 16216 18528
rect 16280 18464 16296 18528
rect 16360 18464 16376 18528
rect 16440 18464 16456 18528
rect 16520 18464 16528 18528
rect 16208 17440 16528 18464
rect 16208 17376 16216 17440
rect 16280 17376 16296 17440
rect 16360 17376 16376 17440
rect 16440 17376 16456 17440
rect 16520 17376 16528 17440
rect 16208 16352 16528 17376
rect 16208 16288 16216 16352
rect 16280 16288 16296 16352
rect 16360 16288 16376 16352
rect 16440 16288 16456 16352
rect 16520 16288 16528 16352
rect 16208 15264 16528 16288
rect 16208 15200 16216 15264
rect 16280 15200 16296 15264
rect 16360 15200 16376 15264
rect 16440 15200 16456 15264
rect 16520 15200 16528 15264
rect 16208 14176 16528 15200
rect 16208 14112 16216 14176
rect 16280 14112 16296 14176
rect 16360 14112 16376 14176
rect 16440 14112 16456 14176
rect 16520 14112 16528 14176
rect 16208 13088 16528 14112
rect 16208 13024 16216 13088
rect 16280 13024 16296 13088
rect 16360 13024 16376 13088
rect 16440 13024 16456 13088
rect 16520 13024 16528 13088
rect 16208 12000 16528 13024
rect 16208 11936 16216 12000
rect 16280 11936 16296 12000
rect 16360 11936 16376 12000
rect 16440 11936 16456 12000
rect 16520 11936 16528 12000
rect 16208 10912 16528 11936
rect 16208 10848 16216 10912
rect 16280 10848 16296 10912
rect 16360 10848 16376 10912
rect 16440 10848 16456 10912
rect 16520 10848 16528 10912
rect 16208 9824 16528 10848
rect 16208 9760 16216 9824
rect 16280 9760 16296 9824
rect 16360 9760 16376 9824
rect 16440 9760 16456 9824
rect 16520 9760 16528 9824
rect 16208 8736 16528 9760
rect 16208 8672 16216 8736
rect 16280 8672 16296 8736
rect 16360 8672 16376 8736
rect 16440 8672 16456 8736
rect 16520 8672 16528 8736
rect 16208 7648 16528 8672
rect 16208 7584 16216 7648
rect 16280 7584 16296 7648
rect 16360 7584 16376 7648
rect 16440 7584 16456 7648
rect 16520 7584 16528 7648
rect 16208 6560 16528 7584
rect 16208 6496 16216 6560
rect 16280 6496 16296 6560
rect 16360 6496 16376 6560
rect 16440 6496 16456 6560
rect 16520 6496 16528 6560
rect 16208 5472 16528 6496
rect 16208 5408 16216 5472
rect 16280 5408 16296 5472
rect 16360 5408 16376 5472
rect 16440 5408 16456 5472
rect 16520 5408 16528 5472
rect 16208 4384 16528 5408
rect 16208 4320 16216 4384
rect 16280 4320 16296 4384
rect 16360 4320 16376 4384
rect 16440 4320 16456 4384
rect 16520 4320 16528 4384
rect 16208 3296 16528 4320
rect 16208 3232 16216 3296
rect 16280 3232 16296 3296
rect 16360 3232 16376 3296
rect 16440 3232 16456 3296
rect 16520 3232 16528 3296
rect 16208 2208 16528 3232
rect 16208 2144 16216 2208
rect 16280 2144 16296 2208
rect 16360 2144 16376 2208
rect 16440 2144 16456 2208
rect 16520 2144 16528 2208
rect 16208 1120 16528 2144
rect 16208 1056 16216 1120
rect 16280 1056 16296 1120
rect 16360 1056 16376 1120
rect 16440 1056 16456 1120
rect 16520 1056 16528 1120
rect 16208 1040 16528 1056
rect 20208 20160 20528 20720
rect 20208 20096 20216 20160
rect 20280 20096 20296 20160
rect 20360 20096 20376 20160
rect 20440 20096 20456 20160
rect 20520 20096 20528 20160
rect 20208 19072 20528 20096
rect 20208 19008 20216 19072
rect 20280 19008 20296 19072
rect 20360 19008 20376 19072
rect 20440 19008 20456 19072
rect 20520 19008 20528 19072
rect 20208 17984 20528 19008
rect 20208 17920 20216 17984
rect 20280 17920 20296 17984
rect 20360 17920 20376 17984
rect 20440 17920 20456 17984
rect 20520 17920 20528 17984
rect 20208 16896 20528 17920
rect 20208 16832 20216 16896
rect 20280 16832 20296 16896
rect 20360 16832 20376 16896
rect 20440 16832 20456 16896
rect 20520 16832 20528 16896
rect 20208 15808 20528 16832
rect 20208 15744 20216 15808
rect 20280 15744 20296 15808
rect 20360 15744 20376 15808
rect 20440 15744 20456 15808
rect 20520 15744 20528 15808
rect 20208 14720 20528 15744
rect 20208 14656 20216 14720
rect 20280 14656 20296 14720
rect 20360 14656 20376 14720
rect 20440 14656 20456 14720
rect 20520 14656 20528 14720
rect 20208 13632 20528 14656
rect 20208 13568 20216 13632
rect 20280 13568 20296 13632
rect 20360 13568 20376 13632
rect 20440 13568 20456 13632
rect 20520 13568 20528 13632
rect 20208 12544 20528 13568
rect 20208 12480 20216 12544
rect 20280 12480 20296 12544
rect 20360 12480 20376 12544
rect 20440 12480 20456 12544
rect 20520 12480 20528 12544
rect 20208 11456 20528 12480
rect 20208 11392 20216 11456
rect 20280 11392 20296 11456
rect 20360 11392 20376 11456
rect 20440 11392 20456 11456
rect 20520 11392 20528 11456
rect 20208 10368 20528 11392
rect 20208 10304 20216 10368
rect 20280 10304 20296 10368
rect 20360 10304 20376 10368
rect 20440 10304 20456 10368
rect 20520 10304 20528 10368
rect 20208 9280 20528 10304
rect 20208 9216 20216 9280
rect 20280 9216 20296 9280
rect 20360 9216 20376 9280
rect 20440 9216 20456 9280
rect 20520 9216 20528 9280
rect 20208 8192 20528 9216
rect 20208 8128 20216 8192
rect 20280 8128 20296 8192
rect 20360 8128 20376 8192
rect 20440 8128 20456 8192
rect 20520 8128 20528 8192
rect 20208 7104 20528 8128
rect 20208 7040 20216 7104
rect 20280 7040 20296 7104
rect 20360 7040 20376 7104
rect 20440 7040 20456 7104
rect 20520 7040 20528 7104
rect 20208 6016 20528 7040
rect 20208 5952 20216 6016
rect 20280 5952 20296 6016
rect 20360 5952 20376 6016
rect 20440 5952 20456 6016
rect 20520 5952 20528 6016
rect 20208 4928 20528 5952
rect 20208 4864 20216 4928
rect 20280 4864 20296 4928
rect 20360 4864 20376 4928
rect 20440 4864 20456 4928
rect 20520 4864 20528 4928
rect 20208 3840 20528 4864
rect 20208 3776 20216 3840
rect 20280 3776 20296 3840
rect 20360 3776 20376 3840
rect 20440 3776 20456 3840
rect 20520 3776 20528 3840
rect 20208 2752 20528 3776
rect 20208 2688 20216 2752
rect 20280 2688 20296 2752
rect 20360 2688 20376 2752
rect 20440 2688 20456 2752
rect 20520 2688 20528 2752
rect 20208 1664 20528 2688
rect 20208 1600 20216 1664
rect 20280 1600 20296 1664
rect 20360 1600 20376 1664
rect 20440 1600 20456 1664
rect 20520 1600 20528 1664
rect 20208 1040 20528 1600
rect 24208 20704 24528 20720
rect 24208 20640 24216 20704
rect 24280 20640 24296 20704
rect 24360 20640 24376 20704
rect 24440 20640 24456 20704
rect 24520 20640 24528 20704
rect 24208 19616 24528 20640
rect 24208 19552 24216 19616
rect 24280 19552 24296 19616
rect 24360 19552 24376 19616
rect 24440 19552 24456 19616
rect 24520 19552 24528 19616
rect 24208 18528 24528 19552
rect 24208 18464 24216 18528
rect 24280 18464 24296 18528
rect 24360 18464 24376 18528
rect 24440 18464 24456 18528
rect 24520 18464 24528 18528
rect 24208 17440 24528 18464
rect 24208 17376 24216 17440
rect 24280 17376 24296 17440
rect 24360 17376 24376 17440
rect 24440 17376 24456 17440
rect 24520 17376 24528 17440
rect 24208 16352 24528 17376
rect 24208 16288 24216 16352
rect 24280 16288 24296 16352
rect 24360 16288 24376 16352
rect 24440 16288 24456 16352
rect 24520 16288 24528 16352
rect 24208 15264 24528 16288
rect 24208 15200 24216 15264
rect 24280 15200 24296 15264
rect 24360 15200 24376 15264
rect 24440 15200 24456 15264
rect 24520 15200 24528 15264
rect 24208 14176 24528 15200
rect 24208 14112 24216 14176
rect 24280 14112 24296 14176
rect 24360 14112 24376 14176
rect 24440 14112 24456 14176
rect 24520 14112 24528 14176
rect 24208 13088 24528 14112
rect 24208 13024 24216 13088
rect 24280 13024 24296 13088
rect 24360 13024 24376 13088
rect 24440 13024 24456 13088
rect 24520 13024 24528 13088
rect 24208 12000 24528 13024
rect 24208 11936 24216 12000
rect 24280 11936 24296 12000
rect 24360 11936 24376 12000
rect 24440 11936 24456 12000
rect 24520 11936 24528 12000
rect 24208 10912 24528 11936
rect 24208 10848 24216 10912
rect 24280 10848 24296 10912
rect 24360 10848 24376 10912
rect 24440 10848 24456 10912
rect 24520 10848 24528 10912
rect 24208 9824 24528 10848
rect 24208 9760 24216 9824
rect 24280 9760 24296 9824
rect 24360 9760 24376 9824
rect 24440 9760 24456 9824
rect 24520 9760 24528 9824
rect 24208 8736 24528 9760
rect 24208 8672 24216 8736
rect 24280 8672 24296 8736
rect 24360 8672 24376 8736
rect 24440 8672 24456 8736
rect 24520 8672 24528 8736
rect 24208 7648 24528 8672
rect 24208 7584 24216 7648
rect 24280 7584 24296 7648
rect 24360 7584 24376 7648
rect 24440 7584 24456 7648
rect 24520 7584 24528 7648
rect 24208 6560 24528 7584
rect 24208 6496 24216 6560
rect 24280 6496 24296 6560
rect 24360 6496 24376 6560
rect 24440 6496 24456 6560
rect 24520 6496 24528 6560
rect 24208 5472 24528 6496
rect 24208 5408 24216 5472
rect 24280 5408 24296 5472
rect 24360 5408 24376 5472
rect 24440 5408 24456 5472
rect 24520 5408 24528 5472
rect 24208 4384 24528 5408
rect 24208 4320 24216 4384
rect 24280 4320 24296 4384
rect 24360 4320 24376 4384
rect 24440 4320 24456 4384
rect 24520 4320 24528 4384
rect 24208 3296 24528 4320
rect 24208 3232 24216 3296
rect 24280 3232 24296 3296
rect 24360 3232 24376 3296
rect 24440 3232 24456 3296
rect 24520 3232 24528 3296
rect 24208 2208 24528 3232
rect 24208 2144 24216 2208
rect 24280 2144 24296 2208
rect 24360 2144 24376 2208
rect 24440 2144 24456 2208
rect 24520 2144 24528 2208
rect 24208 1120 24528 2144
rect 24208 1056 24216 1120
rect 24280 1056 24296 1120
rect 24360 1056 24376 1120
rect 24440 1056 24456 1120
rect 24520 1056 24528 1120
rect 24208 1040 24528 1056
use sky130_fd_sc_hd__nand2b_1  _411_
timestamp -3599
transform -1 0 4416 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _412_
timestamp -3599
transform 1 0 6348 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _413_
timestamp -3599
transform 1 0 5520 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _414_
timestamp -3599
transform 1 0 6992 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _415_
timestamp -3599
transform 1 0 5428 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _416_
timestamp -3599
transform -1 0 6808 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _417_
timestamp -3599
transform -1 0 7728 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _418_
timestamp -3599
transform -1 0 6164 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _419_
timestamp -3599
transform -1 0 4232 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _420_
timestamp -3599
transform 1 0 5244 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _421_
timestamp -3599
transform 1 0 6440 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _422_
timestamp -3599
transform -1 0 6164 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _423_
timestamp -3599
transform 1 0 4416 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _424_
timestamp -3599
transform 1 0 5704 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _425_
timestamp -3599
transform -1 0 8096 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _426_
timestamp -3599
transform 1 0 5980 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _427_
timestamp -3599
transform 1 0 8280 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _428_
timestamp -3599
transform -1 0 6900 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _429_
timestamp -3599
transform -1 0 8924 0 -1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _430_
timestamp -3599
transform -1 0 9568 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _431_
timestamp -3599
transform 1 0 6440 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _432_
timestamp -3599
transform 1 0 7544 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _433_
timestamp -3599
transform -1 0 8188 0 1 1088
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _434_
timestamp -3599
transform 1 0 8372 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _435_
timestamp -3599
transform 1 0 7176 0 -1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _436_
timestamp -3599
transform 1 0 6808 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _437_
timestamp -3599
transform 1 0 8004 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _438_
timestamp -3599
transform 1 0 8372 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _439_
timestamp -3599
transform -1 0 7820 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _440_
timestamp -3599
transform 1 0 8004 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _441_
timestamp -3599
transform 1 0 7360 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _442_
timestamp -3599
transform 1 0 7268 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _443_
timestamp -3599
transform 1 0 7084 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nand2b_1  _444_
timestamp -3599
transform 1 0 5244 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _445_
timestamp -3599
transform 1 0 5244 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _446_
timestamp -3599
transform -1 0 5612 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _447_
timestamp -3599
transform -1 0 5704 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _448_
timestamp -3599
transform 1 0 4416 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _449_
timestamp -3599
transform 1 0 5888 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _450_
timestamp -3599
transform -1 0 6808 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _451_
timestamp -3599
transform 1 0 5520 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _452_
timestamp -3599
transform 1 0 6072 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _453_
timestamp -3599
transform -1 0 6808 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _454_
timestamp -3599
transform -1 0 5244 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _455_
timestamp -3599
transform 1 0 6256 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _456_
timestamp -3599
transform 1 0 4324 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _457_
timestamp -3599
transform 1 0 4784 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _458_
timestamp -3599
transform 1 0 16192 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _459_
timestamp -3599
transform -1 0 17112 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _460_
timestamp -3599
transform -1 0 7636 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _461_
timestamp -3599
transform -1 0 6072 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _462_
timestamp -3599
transform -1 0 5888 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _463_
timestamp -3599
transform -1 0 4140 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _464_
timestamp -3599
transform -1 0 4508 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _465_
timestamp -3599
transform 1 0 2760 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _466_
timestamp -3599
transform 1 0 2208 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _467_
timestamp -3599
transform -1 0 5244 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _468_
timestamp -3599
transform 1 0 2576 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _469_
timestamp -3599
transform 1 0 2024 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _470_
timestamp -3599
transform -1 0 5336 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _471_
timestamp -3599
transform -1 0 5060 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _472_
timestamp -3599
transform 1 0 2576 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _473_
timestamp -3599
transform 1 0 2024 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _474_
timestamp -3599
transform -1 0 4968 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _475_
timestamp -3599
transform 1 0 2760 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _476_
timestamp -3599
transform 1 0 2116 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _477_
timestamp -3599
transform -1 0 6164 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _478_
timestamp -3599
transform -1 0 7084 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _479_
timestamp -3599
transform 1 0 3496 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _480_
timestamp -3599
transform 1 0 2024 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _481_
timestamp -3599
transform -1 0 6348 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _482_
timestamp -3599
transform -1 0 7176 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _483_
timestamp -3599
transform -1 0 8188 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _484_
timestamp -3599
transform 1 0 6440 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _485_
timestamp -3599
transform 1 0 2208 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _486_
timestamp -3599
transform -1 0 6164 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _487_
timestamp -3599
transform -1 0 7360 0 1 1088
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _488_
timestamp -3599
transform 1 0 6348 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _489_
timestamp -3599
transform 1 0 3312 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _490_
timestamp -3599
transform -1 0 16192 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _491_
timestamp -3599
transform 1 0 11316 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _492_
timestamp -3599
transform -1 0 10856 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _493_
timestamp -3599
transform 1 0 7268 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _494_
timestamp -3599
transform 1 0 6440 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _495_
timestamp -3599
transform 1 0 24472 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _496_
timestamp -3599
transform 1 0 23828 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _497_
timestamp -3599
transform 1 0 23368 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _498_
timestamp -3599
transform 1 0 23184 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _499_
timestamp -3599
transform 1 0 20700 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _500_
timestamp -3599
transform -1 0 21068 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _501_
timestamp -3599
transform 1 0 17296 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _502_
timestamp -3599
transform 1 0 16836 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _503_
timestamp -3599
transform -1 0 19228 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _504_
timestamp -3599
transform 1 0 19320 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _505_
timestamp -3599
transform 1 0 14168 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _506_
timestamp -3599
transform -1 0 15272 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _507_
timestamp -3599
transform 1 0 15916 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _508_
timestamp -3599
transform 1 0 12696 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _509_
timestamp -3599
transform -1 0 12512 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _510_
timestamp -3599
transform 1 0 11868 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _511_
timestamp -3599
transform 1 0 11592 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _512_
timestamp -3599
transform 1 0 12236 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _513_
timestamp -3599
transform 1 0 11868 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _514_
timestamp -3599
transform 1 0 12696 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _515_
timestamp -3599
transform 1 0 12236 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _516_
timestamp -3599
transform 1 0 11592 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _517_
timestamp -3599
transform 1 0 11040 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _518_
timestamp -3599
transform 1 0 11868 0 -1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _519_
timestamp -3599
transform 1 0 11592 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _520_
timestamp -3599
transform 1 0 16008 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _521_
timestamp -3599
transform 1 0 23000 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _522_
timestamp -3599
transform -1 0 22816 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _523_
timestamp -3599
transform 1 0 22172 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _524_
timestamp -3599
transform -1 0 21988 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _525_
timestamp -3599
transform 1 0 20516 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _526_
timestamp -3599
transform -1 0 20332 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _527_
timestamp -3599
transform 1 0 16928 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _528_
timestamp -3599
transform -1 0 17020 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _529_
timestamp -3599
transform -1 0 18860 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _530_
timestamp -3599
transform 1 0 18768 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _531_
timestamp -3599
transform 1 0 14904 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _532_
timestamp -3599
transform 1 0 14628 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _533_
timestamp -3599
transform 1 0 23368 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _534_
timestamp -3599
transform -1 0 22356 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _535_
timestamp -3599
transform 1 0 16744 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _536_
timestamp -3599
transform 1 0 21896 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _537_
timestamp -3599
transform 1 0 21344 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _538_
timestamp -3599
transform 1 0 15548 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _539_
timestamp -3599
transform 1 0 15088 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _540_
timestamp -3599
transform 1 0 14628 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _541_
timestamp -3599
transform -1 0 13984 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _542_
timestamp -3599
transform 1 0 17572 0 1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _543_
timestamp -3599
transform 1 0 17020 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _544_
timestamp -3599
transform 1 0 14536 0 1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _545_
timestamp -3599
transform -1 0 14444 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _546_
timestamp -3599
transform 1 0 7728 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _547_
timestamp -3599
transform -1 0 8740 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _548_
timestamp -3599
transform 1 0 7820 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__inv_1  _549_
timestamp -3599
transform 1 0 7360 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _550_
timestamp -3599
transform -1 0 7544 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _551_
timestamp -3599
transform 1 0 7360 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _552_
timestamp -3599
transform -1 0 9016 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _553_
timestamp -3599
transform -1 0 11224 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _554_
timestamp -3599
transform -1 0 9476 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _555_
timestamp -3599
transform -1 0 8740 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _556_
timestamp -3599
transform 1 0 7636 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _557_
timestamp -3599
transform 1 0 10120 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _558_
timestamp -3599
transform 1 0 9200 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _559_
timestamp -3599
transform 1 0 8924 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _560_
timestamp -3599
transform 1 0 9752 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nand3b_1  _561_
timestamp -3599
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _562_
timestamp -3599
transform 1 0 24472 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _563_
timestamp -3599
transform 1 0 24380 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _564_
timestamp -3599
transform 1 0 24472 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _565_
timestamp -3599
transform -1 0 23184 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _566_
timestamp -3599
transform 1 0 20332 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _567_
timestamp -3599
transform 1 0 19872 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _568_
timestamp -3599
transform -1 0 17940 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _569_
timestamp -3599
transform 1 0 17480 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _570_
timestamp -3599
transform 1 0 19320 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _571_
timestamp -3599
transform 1 0 18492 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _572_
timestamp -3599
transform 1 0 14444 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _573_
timestamp -3599
transform 1 0 13616 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _574_
timestamp -3599
transform -1 0 10488 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _575_
timestamp -3599
transform -1 0 10304 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _576_
timestamp -3599
transform 1 0 7912 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _577_
timestamp -3599
transform 1 0 7636 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _578_
timestamp -3599
transform 1 0 10396 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _579_
timestamp -3599
transform 1 0 10212 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _580_
timestamp -3599
transform 1 0 9016 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _581_
timestamp -3599
transform 1 0 8096 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _582_
timestamp -3599
transform 1 0 11592 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _583_
timestamp -3599
transform -1 0 11776 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _584_
timestamp -3599
transform -1 0 10764 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _585_
timestamp -3599
transform 1 0 10488 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _586_
timestamp -3599
transform 1 0 23184 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _587_
timestamp -3599
transform 1 0 22908 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _588_
timestamp -3599
transform 1 0 21896 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _589_
timestamp -3599
transform 1 0 21160 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _590_
timestamp -3599
transform 1 0 16744 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _591_
timestamp -3599
transform 1 0 17848 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _592_
timestamp -3599
transform 1 0 17480 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _593_
timestamp -3599
transform -1 0 17756 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _594_
timestamp -3599
transform 1 0 18216 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _595_
timestamp -3599
transform 1 0 19320 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _596_
timestamp -3599
transform -1 0 19044 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _597_
timestamp -3599
transform 1 0 14720 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _598_
timestamp -3599
transform -1 0 14444 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _599_
timestamp -3599
transform 1 0 19320 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _600_
timestamp -3599
transform -1 0 19780 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _601_
timestamp -3599
transform 1 0 18216 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _602_
timestamp -3599
transform -1 0 18032 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _603_
timestamp -3599
transform 1 0 19780 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _604_
timestamp -3599
transform -1 0 19596 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _605_
timestamp -3599
transform -1 0 16468 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _606_
timestamp -3599
transform 1 0 17204 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _607_
timestamp -3599
transform -1 0 16100 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _608_
timestamp -3599
transform -1 0 17020 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _609_
timestamp -3599
transform 1 0 13616 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _610_
timestamp -3599
transform -1 0 13432 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _611_
timestamp -3599
transform 1 0 3496 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _612_
timestamp -3599
transform 1 0 5060 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _613_
timestamp -3599
transform -1 0 4600 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _614_
timestamp -3599
transform 1 0 3128 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _615_
timestamp -3599
transform -1 0 5888 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _616_
timestamp -3599
transform 1 0 5704 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _617_
timestamp -3599
transform 1 0 3220 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _618_
timestamp -3599
transform 1 0 6164 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand4_1  _619_
timestamp -3599
transform 1 0 6808 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _620_
timestamp -3599
transform 1 0 3864 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _621_
timestamp -3599
transform 1 0 4968 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _622_
timestamp -3599
transform 1 0 4140 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _623_
timestamp -3599
transform 1 0 4968 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__and4bb_1  _624_
timestamp -3599
transform 1 0 3956 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__inv_1  _625_
timestamp -3599
transform 1 0 3956 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _626_
timestamp -3599
transform -1 0 3588 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _627_
timestamp -3599
transform -1 0 4968 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _628_
timestamp -3599
transform -1 0 3588 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _629_
timestamp -3599
transform 1 0 2300 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _630_
timestamp -3599
transform -1 0 5980 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _631_
timestamp -3599
transform -1 0 5060 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _632_
timestamp -3599
transform -1 0 5428 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _633_
timestamp -3599
transform 1 0 3864 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _634_
timestamp -3599
transform 1 0 3680 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _635_
timestamp -3599
transform 1 0 4508 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_2  _636_
timestamp -3599
transform 1 0 3956 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _637_
timestamp -3599
transform 1 0 5520 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _638_
timestamp -3599
transform -1 0 10764 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _639_
timestamp -3599
transform -1 0 8372 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _640_
timestamp -3599
transform -1 0 5336 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _641_
timestamp -3599
transform 1 0 4692 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _642_
timestamp -3599
transform -1 0 4600 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _643_
timestamp -3599
transform -1 0 2484 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _644_
timestamp -3599
transform 1 0 3864 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _645_
timestamp -3599
transform -1 0 4048 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _646_
timestamp -3599
transform -1 0 4784 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _647_
timestamp -3599
transform 1 0 4692 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _648_
timestamp -3599
transform -1 0 6072 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _649_
timestamp -3599
transform 1 0 6440 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _650_
timestamp -3599
transform -1 0 7820 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _651_
timestamp -3599
transform 1 0 10948 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _652_
timestamp -3599
transform 1 0 10948 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nand2b_1  _653_
timestamp -3599
transform -1 0 6072 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _654_
timestamp -3599
transform 1 0 4600 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _655_
timestamp -3599
transform -1 0 5060 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _656_
timestamp -3599
transform 1 0 4876 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _657_
timestamp -3599
transform 1 0 9568 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a41o_1  _658_
timestamp -3599
transform 1 0 9108 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nand2b_1  _659_
timestamp -3599
transform -1 0 8556 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _660_
timestamp -3599
transform 1 0 12236 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2b_1  _661_
timestamp -3599
transform 1 0 13064 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _662_
timestamp -3599
transform 1 0 9844 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _663_
timestamp -3599
transform 1 0 8372 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _664_
timestamp -3599
transform -1 0 5428 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nand3b_1  _665_
timestamp -3599
transform 1 0 5520 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nand3b_2  _666_
timestamp -3599
transform 1 0 6256 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _667_
timestamp -3599
transform -1 0 9660 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _668_
timestamp -3599
transform -1 0 13248 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _669_
timestamp -3599
transform 1 0 11408 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _670_
timestamp -3599
transform 1 0 11684 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _671_
timestamp -3599
transform -1 0 13800 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _672_
timestamp -3599
transform -1 0 14444 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _673_
timestamp -3599
transform -1 0 12144 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _674_
timestamp -3599
transform 1 0 10120 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _675_
timestamp -3599
transform 1 0 10120 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _676_
timestamp -3599
transform -1 0 9476 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _677_
timestamp -3599
transform 1 0 8740 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _678_
timestamp -3599
transform -1 0 7912 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _679_
timestamp -3599
transform 1 0 7084 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _680_
timestamp -3599
transform -1 0 6900 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _681_
timestamp -3599
transform 1 0 6440 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _682_
timestamp -3599
transform 1 0 5520 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _683_
timestamp -3599
transform -1 0 7912 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _684_
timestamp -3599
transform -1 0 8372 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _685_
timestamp -3599
transform -1 0 4508 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _686_
timestamp -3599
transform -1 0 3956 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _687_
timestamp -3599
transform 1 0 2944 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _688_
timestamp -3599
transform 1 0 6072 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _689_
timestamp -3599
transform 1 0 3864 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _690_
timestamp -3599
transform -1 0 3404 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _691_
timestamp -3599
transform 1 0 2944 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _692_
timestamp -3599
transform 1 0 7084 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _693_
timestamp -3599
transform -1 0 7084 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _694_
timestamp -3599
transform 1 0 11040 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _695_
timestamp -3599
transform 1 0 11040 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _696_
timestamp -3599
transform -1 0 13248 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _697_
timestamp -3599
transform -1 0 13892 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _698_
timestamp -3599
transform -1 0 12880 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _699_
timestamp -3599
transform -1 0 13248 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _700_
timestamp -3599
transform 1 0 12788 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _701_
timestamp -3599
transform -1 0 11316 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _702_
timestamp -3599
transform 1 0 10212 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _703_
timestamp -3599
transform -1 0 12236 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _704_
timestamp -3599
transform -1 0 11408 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nand3b_1  _705_
timestamp -3599
transform -1 0 13064 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _706_
timestamp -3599
transform 1 0 11316 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _707_
timestamp -3599
transform -1 0 8648 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _708_
timestamp -3599
transform 1 0 8740 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _709_
timestamp -3599
transform -1 0 7912 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _710_
timestamp -3599
transform -1 0 6164 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _711_
timestamp -3599
transform -1 0 10304 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _712_
timestamp -3599
transform 1 0 10212 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _713_
timestamp -3599
transform 1 0 9660 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _714_
timestamp -3599
transform -1 0 4508 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _715_
timestamp -3599
transform -1 0 4876 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _716_
timestamp -3599
transform 1 0 6440 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _717_
timestamp -3599
transform 1 0 5704 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _718_
timestamp -3599
transform -1 0 5888 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_2  _719_
timestamp -3599
transform -1 0 12512 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _720_
timestamp -3599
transform -1 0 9844 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _721_
timestamp -3599
transform 1 0 8832 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _722_
timestamp -3599
transform -1 0 13800 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _723_
timestamp -3599
transform 1 0 14168 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _724_
timestamp -3599
transform -1 0 14996 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _725_
timestamp -3599
transform -1 0 13800 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _726_
timestamp -3599
transform -1 0 15732 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_2  _727_
timestamp -3599
transform 1 0 14168 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _728_
timestamp -3599
transform 1 0 12696 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _729_
timestamp -3599
transform -1 0 14444 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _730_
timestamp -3599
transform 1 0 13984 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _731_
timestamp -3599
transform 1 0 9016 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _732_
timestamp -3599
transform 1 0 8832 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _733_
timestamp -3599
transform 1 0 10396 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _734_
timestamp -3599
transform -1 0 12604 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _735_
timestamp -3599
transform 1 0 10028 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _736_
timestamp -3599
transform -1 0 11316 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _737_
timestamp -3599
transform -1 0 11132 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _738_
timestamp -3599
transform -1 0 11868 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _739_
timestamp -3599
transform -1 0 10764 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _740_
timestamp -3599
transform -1 0 12328 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _741_
timestamp -3599
transform -1 0 11776 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _742_
timestamp -3599
transform -1 0 10212 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _743_
timestamp -3599
transform 1 0 7912 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _744_
timestamp -3599
transform 1 0 9016 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _745_
timestamp -3599
transform 1 0 8464 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _746_
timestamp -3599
transform 1 0 9660 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _747_
timestamp -3599
transform -1 0 9476 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _748_
timestamp -3599
transform 1 0 9016 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _749_
timestamp -3599
transform -1 0 12328 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _750_
timestamp -3599
transform 1 0 12144 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_1  _751_
timestamp -3599
transform 1 0 11040 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _752_
timestamp -3599
transform -1 0 11316 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nand2b_1  _753_
timestamp -3599
transform -1 0 12880 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _754_
timestamp -3599
transform 1 0 11592 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _755_
timestamp -3599
transform -1 0 11960 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _756_
timestamp -3599
transform -1 0 13156 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _757_
timestamp -3599
transform -1 0 13616 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _758_
timestamp -3599
transform -1 0 12328 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _759_
timestamp -3599
transform 1 0 15916 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _760_
timestamp -3599
transform 1 0 15916 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _761_
timestamp -3599
transform 1 0 14720 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _762_
timestamp -3599
transform 1 0 11040 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _763_
timestamp -3599
transform 1 0 11040 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _764_
timestamp -3599
transform -1 0 4416 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _765_
timestamp -3599
transform -1 0 2760 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _766_
timestamp -3599
transform 1 0 3220 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _767_
timestamp -3599
transform -1 0 9936 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _768_
timestamp -3599
transform 1 0 8004 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _769_
timestamp -3599
transform -1 0 9936 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _770_
timestamp -3599
transform 1 0 11592 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _771_
timestamp -3599
transform 1 0 14628 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _772_
timestamp -3599
transform 1 0 15364 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _773_
timestamp -3599
transform 1 0 14904 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _774_
timestamp -3599
transform 1 0 14812 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _775_
timestamp -3599
transform 1 0 16744 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _776_
timestamp -3599
transform -1 0 17480 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _777_
timestamp -3599
transform -1 0 18952 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _778_
timestamp -3599
transform -1 0 18492 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _779_
timestamp -3599
transform 1 0 14812 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _780_
timestamp -3599
transform -1 0 20608 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _781_
timestamp -3599
transform -1 0 14536 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _782_
timestamp -3599
transform 1 0 20332 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _783_
timestamp -3599
transform 1 0 16192 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _784_
timestamp -3599
transform -1 0 18216 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _785_
timestamp -3599
transform -1 0 21068 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _786_
timestamp -3599
transform 1 0 21252 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _787_
timestamp -3599
transform 1 0 12144 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _788_
timestamp -3599
transform -1 0 12972 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _789_
timestamp -3599
transform 1 0 10672 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _790_
timestamp -3599
transform -1 0 12696 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _791_
timestamp -3599
transform 1 0 9844 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _792_
timestamp -3599
transform 1 0 11040 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _793_
timestamp -3599
transform 1 0 9200 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _794_
timestamp -3599
transform 1 0 11868 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _795_
timestamp -3599
transform -1 0 13064 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _796_
timestamp -3599
transform -1 0 13984 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _797_
timestamp -3599
transform 1 0 20148 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _798_
timestamp -3599
transform 1 0 19320 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _799_
timestamp -3599
transform -1 0 20608 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _800_
timestamp -3599
transform 1 0 23552 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _801_
timestamp -3599
transform 1 0 23644 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _802_
timestamp -3599
transform -1 0 11224 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _803_
timestamp -3599
transform -1 0 10764 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _804_
timestamp -3599
transform 1 0 13248 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _805_
timestamp -3599
transform 1 0 9200 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _806_
timestamp -3599
transform -1 0 10212 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _807_
timestamp -3599
transform 1 0 9200 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _808_
timestamp -3599
transform 1 0 9660 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _809_
timestamp -3599
transform -1 0 14444 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _810_
timestamp -3599
transform -1 0 13892 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _811_
timestamp -3599
transform -1 0 13432 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _812_
timestamp -3599
transform 1 0 14168 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _813_
timestamp -3599
transform -1 0 16100 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _814_
timestamp -3599
transform 1 0 21896 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _815_
timestamp -3599
transform 1 0 21896 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _816_
timestamp -3599
transform 1 0 15456 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _817_
timestamp -3599
transform 1 0 19320 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _818_
timestamp -3599
transform 1 0 17664 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _819_
timestamp -3599
transform -1 0 21252 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _820_
timestamp -3599
transform -1 0 13432 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _821_
timestamp -3599
transform -1 0 22816 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _822_
timestamp -3599
transform 1 0 24472 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _823_
timestamp -3599
transform -1 0 20792 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _824_
timestamp -3599
transform 1 0 21896 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _825_
timestamp -3599
transform 1 0 16468 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _826_
timestamp -3599
transform -1 0 12880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _827_
timestamp -3599
transform 1 0 12880 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _828_
timestamp -3599
transform 1 0 13248 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _829_
timestamp -3599
transform 1 0 12788 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _830_
timestamp -3599
transform 1 0 12328 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _831_
timestamp -3599
transform 1 0 12052 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _832_
timestamp -3599
transform -1 0 12052 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _833_
timestamp -3599
transform 1 0 15364 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _834_
timestamp -3599
transform -1 0 18124 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _835_
timestamp -3599
transform 1 0 18676 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _836_
timestamp -3599
transform 1 0 12972 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _837_
timestamp -3599
transform -1 0 20516 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _838_
timestamp -3599
transform -1 0 22724 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _839_
timestamp -3599
transform 1 0 23368 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _840_
timestamp -3599
transform -1 0 4692 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _841_
timestamp -3599
transform -1 0 3680 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _842_
timestamp -3599
transform 1 0 2760 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _843_
timestamp -3599
transform -1 0 2852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _844_
timestamp -3599
transform -1 0 2760 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _845_
timestamp -3599
transform -1 0 2392 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _846_
timestamp -3599
transform -1 0 2668 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _847_
timestamp -3599
transform -1 0 2760 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _848_
timestamp -3599
transform -1 0 7084 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _849_
timestamp -3599
transform 1 0 3864 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _850_
timestamp -3599
transform 1 0 1656 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _851_
timestamp -3599
transform 1 0 1748 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _852_
timestamp -3599
transform 1 0 8096 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _853_
timestamp -3599
transform 1 0 6808 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _854_
timestamp -3599
transform 1 0 10120 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _855_
timestamp -3599
transform 1 0 14076 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _856_
timestamp -3599
transform 1 0 14168 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _857_
timestamp -3599
transform 1 0 13340 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _858_
timestamp -3599
transform -1 0 17296 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _859_
timestamp -3599
transform -1 0 17572 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _860_
timestamp -3599
transform 1 0 19320 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _861_
timestamp -3599
transform 1 0 17756 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _862_
timestamp -3599
transform 1 0 19504 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _863_
timestamp -3599
transform 1 0 14168 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _864_
timestamp -3599
transform 1 0 18768 0 -1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _865_
timestamp -3599
transform -1 0 18032 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _866_
timestamp -3599
transform 1 0 16928 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _867_
timestamp -3599
transform 1 0 20424 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _868_
timestamp -3599
transform 1 0 22356 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _869_
timestamp -3599
transform 1 0 9292 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _870_
timestamp -3599
transform 1 0 11684 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _871_
timestamp -3599
transform 1 0 7820 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _872_
timestamp -3599
transform 1 0 9660 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _873_
timestamp -3599
transform 1 0 7452 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _874_
timestamp -3599
transform 1 0 10396 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _875_
timestamp -3599
transform 1 0 13156 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _876_
timestamp -3599
transform 1 0 18124 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _877_
timestamp -3599
transform 1 0 17204 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _878_
timestamp -3599
transform 1 0 19504 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _879_
timestamp -3599
transform 1 0 23092 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _880_
timestamp -3599
transform 1 0 23276 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _881_
timestamp -3599
transform 1 0 9016 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _882_
timestamp -3599
transform 1 0 9200 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _883_
timestamp -3599
transform -1 0 9936 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _884_
timestamp -3599
transform 1 0 9016 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _885_
timestamp -3599
transform 1 0 7176 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _886_
timestamp -3599
transform 1 0 7728 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _887_
timestamp -3599
transform -1 0 15364 0 -1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _888_
timestamp -3599
transform 1 0 16744 0 -1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _889_
timestamp -3599
transform -1 0 16008 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _890_
timestamp -3599
transform 1 0 14444 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _891_
timestamp -3599
transform 1 0 20332 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _892_
timestamp -3599
transform -1 0 23184 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _893_
timestamp -3599
transform 1 0 14168 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _894_
timestamp -3599
transform 1 0 17848 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _895_
timestamp -3599
transform 1 0 16744 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _896_
timestamp -3599
transform 1 0 20148 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _897_
timestamp -3599
transform 1 0 21988 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _898_
timestamp -3599
transform 1 0 23000 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _899_
timestamp -3599
transform 1 0 19780 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _900_
timestamp -3599
transform -1 0 22816 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _901_
timestamp -3599
transform 1 0 14628 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _902_
timestamp -3599
transform 1 0 10856 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _903_
timestamp -3599
transform -1 0 11316 0 -1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _904_
timestamp -3599
transform 1 0 11684 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _905_
timestamp -3599
transform 1 0 11592 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _906_
timestamp -3599
transform 1 0 10948 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _907_
timestamp -3599
transform -1 0 13524 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _908_
timestamp -3599
transform -1 0 15824 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _909_
timestamp -3599
transform -1 0 19228 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _910_
timestamp -3599
transform 1 0 16652 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _911_
timestamp -3599
transform -1 0 21804 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _912_
timestamp -3599
transform 1 0 23000 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _913_
timestamp -3599
transform 1 0 23368 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _914_
timestamp -3599
transform 1 0 3864 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _915_
timestamp -3599
transform 1 0 2852 0 -1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _916_
timestamp -3599
transform 1 0 1656 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _917_
timestamp -3599
transform 1 0 1472 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _918_
timestamp -3599
transform 1 0 1472 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _919_
timestamp -3599
transform 1 0 1472 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _920_
timestamp -3599
transform 1 0 1472 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _921_
timestamp -3599
transform 1 0 1656 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _922_
timestamp -3599
transform -1 0 6164 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp -3599
transform -1 0 10856 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp -3599
transform -1 0 6900 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp -3599
transform -1 0 11040 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp -3599
transform 1 0 12512 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp -3599
transform -1 0 15732 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp -3599
transform -1 0 7636 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp -3599
transform -1 0 14536 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clockp_buffer_0
timestamp -3599
transform -1 0 3312 0 1 1088
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_4  clockp_buffer_1
timestamp -3599
transform 1 0 4416 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout104
timestamp -3599
transform 1 0 14168 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  fanout105
timestamp -3599
transform 1 0 13432 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout106
timestamp -3599
transform 1 0 13524 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout107
timestamp -3599
transform 1 0 14628 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout108
timestamp -3599
transform -1 0 13800 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  fanout109
timestamp -3599
transform 1 0 15640 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout110
timestamp -3599
transform 1 0 12512 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout111
timestamp -3599
transform 1 0 9016 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  fanout112
timestamp -3599
transform -1 0 8740 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout113
timestamp -3599
transform -1 0 9936 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout114
timestamp -3599
transform -1 0 10856 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout115
timestamp -3599
transform 1 0 1748 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout116
timestamp -3599
transform 1 0 9384 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  fanout117
timestamp -3599
transform -1 0 10028 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout118
timestamp -3599
transform -1 0 7360 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  fanout119
timestamp -3599
transform -1 0 8004 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout120
timestamp -3599
transform -1 0 15364 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  fanout121
timestamp -3599
transform -1 0 14260 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout122
timestamp -3599
transform -1 0 9844 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  fanout123
timestamp -3599
transform 1 0 8280 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout124
timestamp -3599
transform 1 0 8832 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout125
timestamp -3599
transform 1 0 13432 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout126
timestamp -3599
transform -1 0 13892 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout127
timestamp -3599
transform 1 0 12236 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout128
timestamp -3599
transform 1 0 15180 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  fanout129
timestamp -3599
transform 1 0 15456 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout130
timestamp -3599
transform 1 0 18492 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout131
timestamp -3599
transform 1 0 19136 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout132
timestamp -3599
transform 1 0 20424 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout133
timestamp -3599
transform 1 0 19596 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  fanout134
timestamp -3599
transform -1 0 18584 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout135
timestamp -3599
transform 1 0 10488 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  fanout136
timestamp -3599
transform 1 0 16100 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout137
timestamp -3599
transform 1 0 16560 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  fanout138
timestamp -3599
transform -1 0 18032 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout139
timestamp -3599
transform -1 0 14444 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3
timestamp -3599
transform 1 0 1380 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24
timestamp -3599
transform 1 0 3312 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29
timestamp -3599
transform 1 0 3772 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37
timestamp -3599
transform 1 0 4508 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43
timestamp 1636964856
transform 1 0 5060 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55
timestamp -3599
transform 1 0 6164 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57
timestamp -3599
transform 1 0 6348 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68
timestamp -3599
transform 1 0 7360 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77
timestamp -3599
transform 1 0 8188 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp -3599
transform 1 0 8648 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85
timestamp -3599
transform 1 0 8924 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92
timestamp 1636964856
transform 1 0 9568 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_104
timestamp -3599
transform 1 0 10672 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp -3599
transform 1 0 11316 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113
timestamp -3599
transform 1 0 11500 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117
timestamp 1636964856
transform 1 0 11868 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_129
timestamp -3599
transform 1 0 12972 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp -3599
transform 1 0 13708 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_141
timestamp -3599
transform 1 0 14076 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_145
timestamp -3599
transform 1 0 14444 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_155
timestamp 1636964856
transform 1 0 15364 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp -3599
transform 1 0 16468 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_169
timestamp -3599
transform 1 0 16652 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_176
timestamp -3599
transform 1 0 17296 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_188
timestamp -3599
transform 1 0 18400 0 1 1088
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1636964856
transform 1 0 19228 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1636964856
transform 1 0 20332 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp -3599
transform 1 0 21436 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1636964856
transform 1 0 21804 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1636964856
transform 1 0 22908 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp -3599
transform 1 0 24012 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1636964856
transform 1 0 24380 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_265
timestamp -3599
transform 1 0 25484 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1636964856
transform 1 0 1380 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_15
timestamp -3599
transform 1 0 2484 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_39
timestamp -3599
transform 1 0 4692 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_47
timestamp -3599
transform 1 0 5428 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp -3599
transform 1 0 6072 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_57
timestamp -3599
transform 1 0 6348 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_64
timestamp -3599
transform 1 0 6992 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_73
timestamp -3599
transform 1 0 7820 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_77
timestamp -3599
transform 1 0 8188 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_85
timestamp -3599
transform 1 0 8924 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp -3599
transform 1 0 11316 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_113
timestamp -3599
transform 1 0 11500 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_126
timestamp -3599
transform 1 0 12696 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_131
timestamp -3599
transform 1 0 13156 0 -1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_155
timestamp 1636964856
transform 1 0 15364 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp -3599
transform 1 0 16468 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_169
timestamp -3599
transform 1 0 16652 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_190
timestamp -3599
transform 1 0 18584 0 -1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_212
timestamp 1636964856
transform 1 0 20608 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1636964856
transform 1 0 21804 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1636964856
transform 1 0 22908 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1636964856
transform 1 0 24012 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_261
timestamp -3599
transform 1 0 25116 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_265
timestamp -3599
transform 1 0 25484 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1636964856
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_15
timestamp -3599
transform 1 0 2484 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_23
timestamp -3599
transform 1 0 3220 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp -3599
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_29
timestamp -3599
transform 1 0 3772 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_50
timestamp -3599
transform 1 0 5704 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_55
timestamp -3599
transform 1 0 6164 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_66
timestamp -3599
transform 1 0 7176 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_77
timestamp -3599
transform 1 0 8188 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_82
timestamp -3599
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1636964856
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_97
timestamp -3599
transform 1 0 10028 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_105
timestamp -3599
transform 1 0 10764 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_126
timestamp -3599
transform 1 0 12696 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_130
timestamp -3599
transform 1 0 13064 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_134
timestamp -3599
transform 1 0 13432 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp -3599
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_141
timestamp -3599
transform 1 0 14076 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_162
timestamp -3599
transform 1 0 16008 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_184
timestamp -3599
transform 1 0 18032 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_189
timestamp -3599
transform 1 0 18492 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp -3599
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_197
timestamp -3599
transform 1 0 19228 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_207
timestamp -3599
transform 1 0 20148 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_212
timestamp 1636964856
transform 1 0 20608 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_224
timestamp 1636964856
transform 1 0 21712 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_236
timestamp 1636964856
transform 1 0 22816 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_248
timestamp -3599
transform 1 0 23920 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1636964856
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_265
timestamp -3599
transform 1 0 25484 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1636964856
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_15
timestamp -3599
transform 1 0 2484 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_23
timestamp -3599
transform 1 0 3220 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_28
timestamp -3599
transform 1 0 3680 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_36
timestamp -3599
transform 1 0 4416 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_46
timestamp -3599
transform 1 0 5336 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_53
timestamp -3599
transform 1 0 5980 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_57
timestamp -3599
transform 1 0 6348 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_65
timestamp -3599
transform 1 0 7084 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_73
timestamp -3599
transform 1 0 7820 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_80
timestamp -3599
transform 1 0 8464 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_107
timestamp -3599
transform 1 0 10948 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp -3599
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_113
timestamp -3599
transform 1 0 11500 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_123
timestamp -3599
transform 1 0 12420 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_128
timestamp -3599
transform 1 0 12880 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_136
timestamp -3599
transform 1 0 13616 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_140
timestamp -3599
transform 1 0 13984 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_145
timestamp -3599
transform 1 0 14444 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_156
timestamp -3599
transform 1 0 15456 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp -3599
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_169
timestamp -3599
transform 1 0 16652 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1636964856
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_193
timestamp -3599
transform 1 0 18860 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_201
timestamp -3599
transform 1 0 19596 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp -3599
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_225
timestamp -3599
transform 1 0 21804 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_229
timestamp 1636964856
transform 1 0 22172 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_241
timestamp 1636964856
transform 1 0 23276 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_253
timestamp 1636964856
transform 1 0 24380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_265
timestamp -3599
transform 1 0 25484 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_3
timestamp -3599
transform 1 0 1380 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_11
timestamp -3599
transform 1 0 2116 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_15
timestamp -3599
transform 1 0 2484 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_21
timestamp -3599
transform 1 0 3036 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp -3599
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_29
timestamp -3599
transform 1 0 3772 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_35
timestamp -3599
transform 1 0 4324 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_39
timestamp 1636964856
transform 1 0 4692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_51
timestamp -3599
transform 1 0 5796 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_57
timestamp -3599
transform 1 0 6348 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_66
timestamp -3599
transform 1 0 7176 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_74
timestamp -3599
transform 1 0 7912 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp -3599
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_85
timestamp -3599
transform 1 0 8924 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1636964856
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_124
timestamp -3599
transform 1 0 12512 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_135
timestamp -3599
transform 1 0 13524 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp -3599
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_141
timestamp -3599
transform 1 0 14076 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_145
timestamp 1636964856
transform 1 0 14444 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_157
timestamp -3599
transform 1 0 15548 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_165
timestamp -3599
transform 1 0 16284 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_170
timestamp -3599
transform 1 0 16744 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_174
timestamp -3599
transform 1 0 17112 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp -3599
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_197
timestamp -3599
transform 1 0 19228 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_201
timestamp -3599
transform 1 0 19596 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_209
timestamp -3599
transform 1 0 20332 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_214
timestamp -3599
transform 1 0 20792 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_236
timestamp -3599
transform 1 0 22816 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_247
timestamp -3599
transform 1 0 23828 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp -3599
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1636964856
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_265
timestamp -3599
transform 1 0 25484 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_3
timestamp -3599
transform 1 0 1380 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_26
timestamp -3599
transform 1 0 3496 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_35
timestamp -3599
transform 1 0 4324 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_42
timestamp 1636964856
transform 1 0 4968 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_54
timestamp -3599
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_57
timestamp -3599
transform 1 0 6348 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_67
timestamp -3599
transform 1 0 7268 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_73
timestamp -3599
transform 1 0 7820 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_79
timestamp -3599
transform 1 0 8372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_92
timestamp -3599
transform 1 0 9568 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_100
timestamp -3599
transform 1 0 10304 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_105
timestamp -3599
transform 1 0 10764 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_110
timestamp -3599
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_113
timestamp -3599
transform 1 0 11500 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_135
timestamp -3599
transform 1 0 13524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_141
timestamp -3599
transform 1 0 14076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_145
timestamp -3599
transform 1 0 14444 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp -3599
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_169
timestamp -3599
transform 1 0 16652 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_173
timestamp -3599
transform 1 0 17020 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_183
timestamp -3599
transform 1 0 17940 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_205
timestamp -3599
transform 1 0 19964 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_210
timestamp -3599
transform 1 0 20424 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp -3599
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp -3599
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1636964856
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_237
timestamp -3599
transform 1 0 22908 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_258
timestamp -3599
transform 1 0 24840 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_3
timestamp -3599
transform 1 0 1380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_11
timestamp -3599
transform 1 0 2116 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_18
timestamp -3599
transform 1 0 2760 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp -3599
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp -3599
transform 1 0 3772 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_34
timestamp -3599
transform 1 0 4232 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_43
timestamp -3599
transform 1 0 5060 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_50
timestamp -3599
transform 1 0 5704 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_60
timestamp -3599
transform 1 0 6624 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_69
timestamp -3599
transform 1 0 7452 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_76
timestamp -3599
transform 1 0 8096 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_81
timestamp -3599
transform 1 0 8556 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_85
timestamp -3599
transform 1 0 8924 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_91
timestamp -3599
transform 1 0 9476 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_99
timestamp -3599
transform 1 0 10212 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_106
timestamp -3599
transform 1 0 10856 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_114
timestamp -3599
transform 1 0 11592 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_120
timestamp -3599
transform 1 0 12144 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_125
timestamp -3599
transform 1 0 12604 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_130
timestamp -3599
transform 1 0 13064 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_134
timestamp -3599
transform 1 0 13432 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp -3599
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_141
timestamp -3599
transform 1 0 14076 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_162
timestamp -3599
transform 1 0 16008 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_170
timestamp -3599
transform 1 0 16744 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_181
timestamp -3599
transform 1 0 17756 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_192
timestamp -3599
transform 1 0 18768 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_197
timestamp -3599
transform 1 0 19228 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_207
timestamp -3599
transform 1 0 20148 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_230
timestamp -3599
transform 1 0 22264 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_235
timestamp -3599
transform 1 0 22724 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_240
timestamp -3599
transform 1 0 23184 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp -3599
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_253
timestamp -3599
transform 1 0 24380 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_263
timestamp -3599
transform 1 0 25300 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3
timestamp -3599
transform 1 0 1380 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_24
timestamp -3599
transform 1 0 3312 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_35
timestamp -3599
transform 1 0 4324 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_45
timestamp -3599
transform 1 0 5244 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_49
timestamp -3599
transform 1 0 5612 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp -3599
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_57
timestamp -3599
transform 1 0 6348 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_65
timestamp -3599
transform 1 0 7084 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_71
timestamp -3599
transform 1 0 7636 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_75
timestamp -3599
transform 1 0 8004 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_96
timestamp -3599
transform 1 0 9936 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_101
timestamp -3599
transform 1 0 10396 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_109
timestamp -3599
transform 1 0 11132 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_113
timestamp -3599
transform 1 0 11500 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_134
timestamp -3599
transform 1 0 13432 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_140
timestamp -3599
transform 1 0 13984 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_146
timestamp -3599
transform 1 0 14536 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_157
timestamp -3599
transform 1 0 15548 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_164
timestamp -3599
transform 1 0 16192 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_169
timestamp -3599
transform 1 0 16652 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_174
timestamp -3599
transform 1 0 17112 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_191
timestamp -3599
transform 1 0 18676 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_195
timestamp -3599
transform 1 0 19044 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_206
timestamp -3599
transform 1 0 20056 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_7_212
timestamp -3599
transform 1 0 20608 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_7_221
timestamp -3599
transform 1 0 21436 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_225
timestamp -3599
transform 1 0 21804 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_235
timestamp -3599
transform 1 0 22724 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_259
timestamp -3599
transform 1 0 24932 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_265
timestamp -3599
transform 1 0 25484 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3
timestamp -3599
transform 1 0 1380 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_9
timestamp -3599
transform 1 0 1932 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_13
timestamp -3599
transform 1 0 2300 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_19
timestamp -3599
transform 1 0 2852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp -3599
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_29
timestamp -3599
transform 1 0 3772 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_35
timestamp -3599
transform 1 0 4324 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_43
timestamp -3599
transform 1 0 5060 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_48
timestamp -3599
transform 1 0 5520 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_57
timestamp -3599
transform 1 0 6348 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_63
timestamp -3599
transform 1 0 6900 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_69
timestamp -3599
transform 1 0 7452 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_75
timestamp -3599
transform 1 0 8004 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp -3599
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_85
timestamp -3599
transform 1 0 8924 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_107
timestamp -3599
transform 1 0 10948 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_115
timestamp -3599
transform 1 0 11684 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_8_130
timestamp -3599
transform 1 0 13064 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_136
timestamp -3599
transform 1 0 13616 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_141
timestamp -3599
transform 1 0 14076 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_149
timestamp -3599
transform 1 0 14812 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_155
timestamp -3599
transform 1 0 15364 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_166
timestamp -3599
transform 1 0 16376 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_192
timestamp -3599
transform 1 0 18768 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_8_197
timestamp -3599
transform 1 0 19228 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_220
timestamp 1636964856
transform 1 0 21344 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_232
timestamp -3599
transform 1 0 22448 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_243
timestamp -3599
transform 1 0 23460 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_248
timestamp -3599
transform 1 0 23920 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1636964856
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_265
timestamp -3599
transform 1 0 25484 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_3
timestamp -3599
transform 1 0 1380 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_14
timestamp -3599
transform 1 0 2392 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_27
timestamp -3599
transform 1 0 3588 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_42
timestamp -3599
transform 1 0 4968 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_50
timestamp -3599
transform 1 0 5704 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp -3599
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_57
timestamp -3599
transform 1 0 6348 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_62
timestamp -3599
transform 1 0 6808 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_70
timestamp -3599
transform 1 0 7544 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_77
timestamp -3599
transform 1 0 8188 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_86
timestamp -3599
transform 1 0 9016 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_94
timestamp -3599
transform 1 0 9752 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_99
timestamp -3599
transform 1 0 10212 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_105
timestamp -3599
transform 1 0 10764 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_110
timestamp -3599
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_113
timestamp -3599
transform 1 0 11500 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_126
timestamp -3599
transform 1 0 12696 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_9_136
timestamp -3599
transform 1 0 13616 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_144
timestamp -3599
transform 1 0 14352 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_165
timestamp -3599
transform 1 0 16284 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_169
timestamp -3599
transform 1 0 16652 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_174
timestamp -3599
transform 1 0 17112 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_181
timestamp -3599
transform 1 0 17756 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_186
timestamp -3599
transform 1 0 18216 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_193
timestamp -3599
transform 1 0 18860 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_201
timestamp -3599
transform 1 0 19596 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_207
timestamp -3599
transform 1 0 20148 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_218
timestamp -3599
transform 1 0 21160 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp -3599
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_225
timestamp -3599
transform 1 0 21804 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_235
timestamp -3599
transform 1 0 22724 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_261
timestamp -3599
transform 1 0 25116 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_265
timestamp -3599
transform 1 0 25484 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_3
timestamp -3599
transform 1 0 1380 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_24
timestamp -3599
transform 1 0 3312 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_29
timestamp -3599
transform 1 0 3772 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_35
timestamp -3599
transform 1 0 4324 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_40
timestamp -3599
transform 1 0 4784 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_49
timestamp -3599
transform 1 0 5612 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_55
timestamp 1636964856
transform 1 0 6164 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_67
timestamp -3599
transform 1 0 7268 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_76
timestamp -3599
transform 1 0 8096 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp -3599
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_85
timestamp -3599
transform 1 0 8924 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_91
timestamp -3599
transform 1 0 9476 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_96
timestamp -3599
transform 1 0 9936 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_104
timestamp -3599
transform 1 0 10672 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_127
timestamp -3599
transform 1 0 12788 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_133
timestamp -3599
transform 1 0 13340 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp -3599
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_141
timestamp -3599
transform 1 0 14076 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_154
timestamp -3599
transform 1 0 15272 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_159
timestamp 1636964856
transform 1 0 15732 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_171
timestamp -3599
transform 1 0 16836 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_179
timestamp -3599
transform 1 0 17572 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_185
timestamp -3599
transform 1 0 18124 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_190
timestamp -3599
transform 1 0 18584 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1636964856
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_229
timestamp -3599
transform 1 0 22172 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_237
timestamp -3599
transform 1 0 22908 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_249
timestamp -3599
transform 1 0 24012 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_253
timestamp -3599
transform 1 0 24380 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_263
timestamp -3599
transform 1 0 25300 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1636964856
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_18
timestamp -3599
transform 1 0 2760 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_26
timestamp -3599
transform 1 0 3496 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_34
timestamp -3599
transform 1 0 4232 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_43
timestamp -3599
transform 1 0 5060 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_52
timestamp -3599
transform 1 0 5888 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_57
timestamp -3599
transform 1 0 6348 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_61
timestamp -3599
transform 1 0 6716 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_70
timestamp -3599
transform 1 0 7544 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_92
timestamp -3599
transform 1 0 9568 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_97
timestamp 1636964856
transform 1 0 10028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_109
timestamp -3599
transform 1 0 11132 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_113
timestamp -3599
transform 1 0 11500 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_117
timestamp -3599
transform 1 0 11868 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_122
timestamp -3599
transform 1 0 12328 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_130
timestamp -3599
transform 1 0 13064 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_151
timestamp -3599
transform 1 0 14996 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_163
timestamp -3599
transform 1 0 16100 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp -3599
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_169
timestamp -3599
transform 1 0 16652 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_174
timestamp -3599
transform 1 0 17112 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_197
timestamp -3599
transform 1 0 19228 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_11_205
timestamp -3599
transform 1 0 19964 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_211
timestamp -3599
transform 1 0 20516 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_222
timestamp -3599
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_225
timestamp -3599
transform 1 0 21804 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_229
timestamp -3599
transform 1 0 22172 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_251
timestamp -3599
transform 1 0 24196 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_256
timestamp -3599
transform 1 0 24656 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_264
timestamp -3599
transform 1 0 25392 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_3
timestamp -3599
transform 1 0 1380 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_14
timestamp -3599
transform 1 0 2392 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_25
timestamp -3599
transform 1 0 3404 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp -3599
transform 1 0 3772 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_38
timestamp -3599
transform 1 0 4600 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_46
timestamp -3599
transform 1 0 5336 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_52
timestamp -3599
transform 1 0 5888 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_58
timestamp -3599
transform 1 0 6440 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_66
timestamp -3599
transform 1 0 7176 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_71
timestamp -3599
transform 1 0 7636 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_79
timestamp -3599
transform 1 0 8372 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp -3599
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_85
timestamp -3599
transform 1 0 8924 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_89
timestamp -3599
transform 1 0 9292 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_94
timestamp -3599
transform 1 0 9752 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_105
timestamp 1636964856
transform 1 0 10764 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_117
timestamp -3599
transform 1 0 11868 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_125
timestamp -3599
transform 1 0 12604 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_130
timestamp -3599
transform 1 0 13064 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp -3599
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_141
timestamp -3599
transform 1 0 14076 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_146
timestamp -3599
transform 1 0 14536 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_153
timestamp -3599
transform 1 0 15180 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_158
timestamp -3599
transform 1 0 15640 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_163
timestamp -3599
transform 1 0 16100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_189
timestamp -3599
transform 1 0 18492 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp -3599
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_197
timestamp -3599
transform 1 0 19228 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_201
timestamp -3599
transform 1 0 19596 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_225
timestamp 1636964856
transform 1 0 21804 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_240
timestamp -3599
transform 1 0 23184 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_245
timestamp -3599
transform 1 0 23644 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_250
timestamp -3599
transform 1 0 24104 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_253
timestamp -3599
transform 1 0 24380 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_263
timestamp -3599
transform 1 0 25300 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_3
timestamp -3599
transform 1 0 1380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_24
timestamp -3599
transform 1 0 3312 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_29
timestamp -3599
transform 1 0 3772 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_40
timestamp -3599
transform 1 0 4784 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_46
timestamp -3599
transform 1 0 5336 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp -3599
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_57
timestamp -3599
transform 1 0 6348 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_65
timestamp -3599
transform 1 0 7084 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_86
timestamp -3599
transform 1 0 9016 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_91
timestamp -3599
transform 1 0 9476 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_102
timestamp -3599
transform 1 0 10488 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_107
timestamp -3599
transform 1 0 10948 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp -3599
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_113
timestamp -3599
transform 1 0 11500 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_119
timestamp -3599
transform 1 0 12052 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_124
timestamp -3599
transform 1 0 12512 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_135
timestamp -3599
transform 1 0 13524 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_139
timestamp -3599
transform 1 0 13892 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_160
timestamp -3599
transform 1 0 15824 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp -3599
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_174
timestamp -3599
transform 1 0 17112 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_185
timestamp -3599
transform 1 0 18124 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_197
timestamp -3599
transform 1 0 19228 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_13_203
timestamp -3599
transform 1 0 19780 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_212
timestamp -3599
transform 1 0 20608 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_217
timestamp -3599
transform 1 0 21068 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_222
timestamp -3599
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_225
timestamp -3599
transform 1 0 21804 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_229
timestamp 1636964856
transform 1 0 22172 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_241
timestamp -3599
transform 1 0 23276 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_262
timestamp -3599
transform 1 0 25208 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_3
timestamp -3599
transform 1 0 1380 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_9
timestamp -3599
transform 1 0 1932 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_13
timestamp -3599
transform 1 0 2300 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_21
timestamp -3599
transform 1 0 3036 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp -3599
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp -3599
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_41
timestamp -3599
transform 1 0 4876 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_46
timestamp -3599
transform 1 0 5336 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_55
timestamp -3599
transform 1 0 6164 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_62
timestamp -3599
transform 1 0 6808 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_67
timestamp -3599
transform 1 0 7268 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp -3599
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp -3599
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_85
timestamp -3599
transform 1 0 8924 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_109
timestamp -3599
transform 1 0 11132 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_135
timestamp -3599
transform 1 0 13524 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp -3599
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_141
timestamp -3599
transform 1 0 14076 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_154
timestamp -3599
transform 1 0 15272 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_159
timestamp -3599
transform 1 0 15732 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_164
timestamp 1636964856
transform 1 0 16192 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_176
timestamp -3599
transform 1 0 17296 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_183
timestamp 1636964856
transform 1 0 17940 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp -3599
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_197
timestamp -3599
transform 1 0 19228 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_207
timestamp -3599
transform 1 0 20148 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_14_214
timestamp -3599
transform 1 0 20792 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_240
timestamp -3599
transform 1 0 23184 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp -3599
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_253
timestamp -3599
transform 1 0 24380 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_257
timestamp -3599
transform 1 0 24748 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_265
timestamp -3599
transform 1 0 25484 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_3
timestamp -3599
transform 1 0 1380 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_9
timestamp -3599
transform 1 0 1932 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_13
timestamp -3599
transform 1 0 2300 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_25
timestamp -3599
transform 1 0 3404 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_40
timestamp -3599
transform 1 0 4784 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_48
timestamp -3599
transform 1 0 5520 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp -3599
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_57
timestamp -3599
transform 1 0 6348 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_62
timestamp -3599
transform 1 0 6808 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_68
timestamp -3599
transform 1 0 7360 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_89
timestamp -3599
transform 1 0 9292 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_100
timestamp -3599
transform 1 0 10304 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_105
timestamp -3599
transform 1 0 10764 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp -3599
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_113
timestamp -3599
transform 1 0 11500 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_120
timestamp 1636964856
transform 1 0 12144 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_132
timestamp -3599
transform 1 0 13248 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_140
timestamp -3599
transform 1 0 13984 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_162
timestamp -3599
transform 1 0 16008 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_169
timestamp -3599
transform 1 0 16652 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_190
timestamp -3599
transform 1 0 18584 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_195
timestamp -3599
transform 1 0 19044 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_199
timestamp -3599
transform 1 0 19412 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_220
timestamp -3599
transform 1 0 21344 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_225
timestamp -3599
transform 1 0 21804 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_231
timestamp -3599
transform 1 0 22356 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_236
timestamp -3599
transform 1 0 22816 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_258
timestamp -3599
transform 1 0 24840 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_3
timestamp -3599
transform 1 0 1380 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_24
timestamp -3599
transform 1 0 3312 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_29
timestamp -3599
transform 1 0 3772 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_36
timestamp -3599
transform 1 0 4416 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_45
timestamp -3599
transform 1 0 5244 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_53
timestamp -3599
transform 1 0 5980 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_60
timestamp -3599
transform 1 0 6624 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_67
timestamp -3599
transform 1 0 7268 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_72
timestamp -3599
transform 1 0 7728 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp -3599
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_85
timestamp -3599
transform 1 0 8924 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_95
timestamp -3599
transform 1 0 9844 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_121
timestamp -3599
transform 1 0 12236 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_126
timestamp -3599
transform 1 0 12696 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_134
timestamp -3599
transform 1 0 13432 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_141
timestamp -3599
transform 1 0 14076 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_146
timestamp -3599
transform 1 0 14536 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_159
timestamp -3599
transform 1 0 15732 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_166
timestamp -3599
transform 1 0 16376 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_16_181
timestamp -3599
transform 1 0 17756 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_193
timestamp -3599
transform 1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_197
timestamp -3599
transform 1 0 19228 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_201
timestamp -3599
transform 1 0 19596 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_16_227
timestamp -3599
transform 1 0 21988 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_236
timestamp -3599
transform 1 0 22816 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_247
timestamp -3599
transform 1 0 23828 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp -3599
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1636964856
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_265
timestamp -3599
transform 1 0 25484 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_3
timestamp -3599
transform 1 0 1380 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_11
timestamp -3599
transform 1 0 2116 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_17_17
timestamp -3599
transform 1 0 2668 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_28
timestamp -3599
transform 1 0 3680 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_37
timestamp -3599
transform 1 0 4508 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_45
timestamp -3599
transform 1 0 5244 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_52
timestamp -3599
transform 1 0 5888 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_57
timestamp -3599
transform 1 0 6348 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_62
timestamp -3599
transform 1 0 6808 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_66
timestamp -3599
transform 1 0 7176 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_71
timestamp -3599
transform 1 0 7636 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_93
timestamp -3599
transform 1 0 9660 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_98
timestamp -3599
transform 1 0 10120 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp -3599
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_113
timestamp -3599
transform 1 0 11500 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_123
timestamp -3599
transform 1 0 12420 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_129
timestamp -3599
transform 1 0 12972 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_134
timestamp -3599
transform 1 0 13432 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_145
timestamp -3599
transform 1 0 14444 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_150
timestamp -3599
transform 1 0 14904 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_163
timestamp -3599
transform 1 0 16100 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp -3599
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_169
timestamp -3599
transform 1 0 16652 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_173
timestamp -3599
transform 1 0 17020 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_181
timestamp -3599
transform 1 0 17756 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_202
timestamp 1636964856
transform 1 0 19688 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_214
timestamp -3599
transform 1 0 20792 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_219
timestamp -3599
transform 1 0 21252 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp -3599
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_225
timestamp -3599
transform 1 0 21804 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_247
timestamp 1636964856
transform 1 0 23828 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_259
timestamp -3599
transform 1 0 24932 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_265
timestamp -3599
transform 1 0 25484 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_3
timestamp -3599
transform 1 0 1380 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_11
timestamp -3599
transform 1 0 2116 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_15
timestamp -3599
transform 1 0 2484 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp -3599
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_29
timestamp -3599
transform 1 0 3772 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_18_42
timestamp -3599
transform 1 0 4968 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_54
timestamp -3599
transform 1 0 6072 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_60
timestamp -3599
transform 1 0 6624 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_65
timestamp -3599
transform 1 0 7084 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_18_74
timestamp -3599
transform 1 0 7912 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_79
timestamp -3599
transform 1 0 8372 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp -3599
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_85
timestamp -3599
transform 1 0 8924 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_91
timestamp -3599
transform 1 0 9476 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_113
timestamp -3599
transform 1 0 11500 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_135
timestamp -3599
transform 1 0 13524 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp -3599
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_141
timestamp -3599
transform 1 0 14076 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_145
timestamp -3599
transform 1 0 14444 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_151
timestamp -3599
transform 1 0 14996 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_155
timestamp -3599
transform 1 0 15364 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_176
timestamp -3599
transform 1 0 17296 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_180
timestamp -3599
transform 1 0 17664 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_184
timestamp -3599
transform 1 0 18032 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp -3599
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_197
timestamp -3599
transform 1 0 19228 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_201
timestamp -3599
transform 1 0 19596 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_205
timestamp -3599
transform 1 0 19964 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_209
timestamp -3599
transform 1 0 20332 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_220
timestamp -3599
transform 1 0 21344 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_227
timestamp -3599
transform 1 0 21988 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_238
timestamp 1636964856
transform 1 0 23000 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_250
timestamp -3599
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1636964856
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_265
timestamp -3599
transform 1 0 25484 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_3
timestamp -3599
transform 1 0 1380 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_26
timestamp -3599
transform 1 0 3496 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_33
timestamp -3599
transform 1 0 4140 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp -3599
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1636964856
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_69
timestamp -3599
transform 1 0 7452 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_75
timestamp -3599
transform 1 0 8004 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_96
timestamp -3599
transform 1 0 9936 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_102
timestamp -3599
transform 1 0 10488 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_106
timestamp -3599
transform 1 0 10856 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp -3599
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_113
timestamp -3599
transform 1 0 11500 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_118
timestamp -3599
transform 1 0 11960 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_124
timestamp -3599
transform 1 0 12512 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_132
timestamp -3599
transform 1 0 13248 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_153
timestamp -3599
transform 1 0 15180 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_157
timestamp -3599
transform 1 0 15548 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp -3599
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_169
timestamp -3599
transform 1 0 16652 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_173
timestamp -3599
transform 1 0 17020 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_178
timestamp -3599
transform 1 0 17480 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_201
timestamp -3599
transform 1 0 19596 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_212
timestamp 1636964856
transform 1 0 20608 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1636964856
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_237
timestamp 1636964856
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_249
timestamp 1636964856
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_261
timestamp -3599
transform 1 0 25116 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_265
timestamp -3599
transform 1 0 25484 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1636964856
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_18
timestamp -3599
transform 1 0 2760 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_26
timestamp -3599
transform 1 0 3496 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp -3599
transform 1 0 3772 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_36
timestamp -3599
transform 1 0 4416 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_47
timestamp -3599
transform 1 0 5428 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_52
timestamp 1636964856
transform 1 0 5888 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_64
timestamp 1636964856
transform 1 0 6992 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_76
timestamp -3599
transform 1 0 8096 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_85
timestamp -3599
transform 1 0 8924 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_20_96
timestamp -3599
transform 1 0 9936 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_106
timestamp -3599
transform 1 0 10856 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_111
timestamp -3599
transform 1 0 11316 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_116
timestamp 1636964856
transform 1 0 11776 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_128
timestamp -3599
transform 1 0 12880 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_20_137
timestamp -3599
transform 1 0 13708 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_141
timestamp -3599
transform 1 0 14076 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_20_152
timestamp -3599
transform 1 0 15088 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_158
timestamp -3599
transform 1 0 15640 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_179
timestamp -3599
transform 1 0 17572 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_184
timestamp -3599
transform 1 0 18032 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_189
timestamp -3599
transform 1 0 18492 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp -3599
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_197
timestamp -3599
transform 1 0 19228 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_218
timestamp 1636964856
transform 1 0 21160 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_230
timestamp 1636964856
transform 1 0 22264 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_242
timestamp -3599
transform 1 0 23368 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_250
timestamp -3599
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1636964856
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_265
timestamp -3599
transform 1 0 25484 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1636964856
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1636964856
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_27
timestamp -3599
transform 1 0 3588 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_32
timestamp -3599
transform 1 0 4048 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_40
timestamp -3599
transform 1 0 4784 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_46
timestamp -3599
transform 1 0 5336 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp -3599
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_57
timestamp -3599
transform 1 0 6348 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_61
timestamp -3599
transform 1 0 6716 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_74
timestamp -3599
transform 1 0 7912 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_79
timestamp -3599
transform 1 0 8372 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_83
timestamp -3599
transform 1 0 8740 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_87
timestamp -3599
transform 1 0 9108 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_91
timestamp -3599
transform 1 0 9476 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_96
timestamp -3599
transform 1 0 9936 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_107
timestamp -3599
transform 1 0 10948 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp -3599
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_113
timestamp -3599
transform 1 0 11500 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_120
timestamp 1636964856
transform 1 0 12144 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_132
timestamp 1636964856
transform 1 0 13248 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_144
timestamp -3599
transform 1 0 14352 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_153
timestamp -3599
transform 1 0 15180 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_158
timestamp -3599
transform 1 0 15640 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp -3599
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_169
timestamp -3599
transform 1 0 16652 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_173
timestamp -3599
transform 1 0 17020 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_178
timestamp 1636964856
transform 1 0 17480 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_190
timestamp 1636964856
transform 1 0 18584 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_202
timestamp 1636964856
transform 1 0 19688 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_214
timestamp -3599
transform 1 0 20792 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp -3599
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_225
timestamp 1636964856
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_237
timestamp 1636964856
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_249
timestamp 1636964856
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_261
timestamp -3599
transform 1 0 25116 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_265
timestamp -3599
transform 1 0 25484 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1636964856
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_15
timestamp -3599
transform 1 0 2484 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_19
timestamp -3599
transform 1 0 2852 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp -3599
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_29
timestamp -3599
transform 1 0 3772 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_37
timestamp -3599
transform 1 0 4508 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_44
timestamp -3599
transform 1 0 5152 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_54
timestamp -3599
transform 1 0 6072 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_65
timestamp -3599
transform 1 0 7084 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_74
timestamp -3599
transform 1 0 7912 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_79
timestamp -3599
transform 1 0 8372 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp -3599
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_85
timestamp -3599
transform 1 0 8924 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_91
timestamp -3599
transform 1 0 9476 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_96
timestamp -3599
transform 1 0 9936 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_118
timestamp -3599
transform 1 0 11960 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_126
timestamp -3599
transform 1 0 12696 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp -3599
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_141
timestamp -3599
transform 1 0 14076 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_162
timestamp -3599
transform 1 0 16008 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_22_172
timestamp 1636964856
transform 1 0 16928 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_184
timestamp 1636964856
transform 1 0 18032 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1636964856
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1636964856
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_221
timestamp 1636964856
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_233
timestamp 1636964856
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp -3599
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp -3599
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1636964856
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_265
timestamp -3599
transform 1 0 25484 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_3
timestamp -3599
transform 1 0 1380 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_15
timestamp -3599
transform 1 0 2484 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_25
timestamp -3599
transform 1 0 3404 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_29
timestamp -3599
transform 1 0 3772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_37
timestamp -3599
transform 1 0 4508 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_46
timestamp -3599
transform 1 0 5336 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp -3599
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_57
timestamp -3599
transform 1 0 6348 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_63
timestamp -3599
transform 1 0 6900 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_74
timestamp -3599
transform 1 0 7912 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_81
timestamp -3599
transform 1 0 8556 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_86
timestamp -3599
transform 1 0 9016 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_93
timestamp -3599
transform 1 0 9660 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_97
timestamp -3599
transform 1 0 10028 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_105
timestamp -3599
transform 1 0 10764 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp -3599
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_113
timestamp -3599
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_122
timestamp -3599
transform 1 0 12328 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_134
timestamp -3599
transform 1 0 13432 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_140
timestamp -3599
transform 1 0 13984 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_161
timestamp -3599
transform 1 0 15916 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp -3599
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1636964856
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1636964856
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_193
timestamp 1636964856
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_205
timestamp 1636964856
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp -3599
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp -3599
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_225
timestamp 1636964856
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_237
timestamp 1636964856
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_249
timestamp 1636964856
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_261
timestamp -3599
transform 1 0 25116 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_265
timestamp -3599
transform 1 0 25484 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_3
timestamp -3599
transform 1 0 1380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp -3599
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_29
timestamp -3599
transform 1 0 3772 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_37
timestamp -3599
transform 1 0 4508 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_46
timestamp -3599
transform 1 0 5336 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_52
timestamp -3599
transform 1 0 5888 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_57
timestamp -3599
transform 1 0 6348 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_63
timestamp -3599
transform 1 0 6900 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_73
timestamp -3599
transform 1 0 7820 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_77
timestamp -3599
transform 1 0 8188 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_81
timestamp -3599
transform 1 0 8556 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_85
timestamp -3599
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_95
timestamp -3599
transform 1 0 9844 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_101
timestamp -3599
transform 1 0 10396 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_105
timestamp -3599
transform 1 0 10764 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_110
timestamp -3599
transform 1 0 11224 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_119
timestamp -3599
transform 1 0 12052 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_132
timestamp -3599
transform 1 0 13248 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp -3599
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_141
timestamp -3599
transform 1 0 14076 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_145
timestamp -3599
transform 1 0 14444 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_150
timestamp -3599
transform 1 0 14904 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_161
timestamp -3599
transform 1 0 15916 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_166
timestamp -3599
transform 1 0 16376 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_173
timestamp 1636964856
transform 1 0 17020 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_185
timestamp -3599
transform 1 0 18124 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_193
timestamp -3599
transform 1 0 18860 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1636964856
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_209
timestamp 1636964856
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_221
timestamp 1636964856
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_233
timestamp 1636964856
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp -3599
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp -3599
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1636964856
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_265
timestamp -3599
transform 1 0 25484 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_3
timestamp -3599
transform 1 0 1380 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_26
timestamp -3599
transform 1 0 3496 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_31
timestamp -3599
transform 1 0 3956 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_38
timestamp -3599
transform 1 0 4600 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_42
timestamp -3599
transform 1 0 4968 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_47
timestamp -3599
transform 1 0 5428 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp -3599
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_57
timestamp -3599
transform 1 0 6348 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_61
timestamp -3599
transform 1 0 6716 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_82
timestamp -3599
transform 1 0 8648 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_95
timestamp -3599
transform 1 0 9844 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_100
timestamp -3599
transform 1 0 10304 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp -3599
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_113
timestamp -3599
transform 1 0 11500 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_117
timestamp -3599
transform 1 0 11868 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_124
timestamp -3599
transform 1 0 12512 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_129
timestamp -3599
transform 1 0 12972 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_25_138
timestamp 1636964856
transform 1 0 13800 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_150
timestamp -3599
transform 1 0 14904 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp -3599
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_169
timestamp -3599
transform 1 0 16652 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_183
timestamp 1636964856
transform 1 0 17940 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_195
timestamp 1636964856
transform 1 0 19044 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_207
timestamp 1636964856
transform 1 0 20148 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_219
timestamp -3599
transform 1 0 21252 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp -3599
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1636964856
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_237
timestamp 1636964856
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_249
timestamp 1636964856
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_261
timestamp -3599
transform 1 0 25116 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_265
timestamp -3599
transform 1 0 25484 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1636964856
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_18
timestamp -3599
transform 1 0 2760 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp -3599
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_29
timestamp -3599
transform 1 0 3772 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_50
timestamp -3599
transform 1 0 5704 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_56
timestamp -3599
transform 1 0 6256 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_60
timestamp -3599
transform 1 0 6624 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_68
timestamp -3599
transform 1 0 7360 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_74
timestamp -3599
transform 1 0 7912 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_78
timestamp -3599
transform 1 0 8280 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp -3599
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_85
timestamp -3599
transform 1 0 8924 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_90
timestamp -3599
transform 1 0 9384 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_97
timestamp -3599
transform 1 0 10028 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_105
timestamp -3599
transform 1 0 10764 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_113
timestamp -3599
transform 1 0 11500 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_124
timestamp -3599
transform 1 0 12512 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_132
timestamp -3599
transform 1 0 13248 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_137
timestamp -3599
transform 1 0 13708 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_141
timestamp -3599
transform 1 0 14076 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_152
timestamp -3599
transform 1 0 15088 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_156
timestamp -3599
transform 1 0 15456 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_168
timestamp 1636964856
transform 1 0 16560 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_180
timestamp 1636964856
transform 1 0 17664 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_192
timestamp -3599
transform 1 0 18768 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1636964856
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_209
timestamp 1636964856
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_221
timestamp 1636964856
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_233
timestamp 1636964856
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp -3599
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp -3599
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1636964856
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_265
timestamp -3599
transform 1 0 25484 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1636964856
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_15
timestamp -3599
transform 1 0 2484 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_27_26
timestamp -3599
transform 1 0 3496 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_32
timestamp -3599
transform 1 0 4048 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_36
timestamp 1636964856
transform 1 0 4416 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_48
timestamp -3599
transform 1 0 5520 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp -3599
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_57
timestamp -3599
transform 1 0 6348 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_63
timestamp -3599
transform 1 0 6900 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_68
timestamp -3599
transform 1 0 7360 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_75
timestamp -3599
transform 1 0 8004 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_91
timestamp -3599
transform 1 0 9476 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_100
timestamp -3599
transform 1 0 10304 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp -3599
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_113
timestamp -3599
transform 1 0 11500 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_121
timestamp -3599
transform 1 0 12236 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_131
timestamp -3599
transform 1 0 13156 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_139
timestamp -3599
transform 1 0 13892 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_145
timestamp -3599
transform 1 0 14444 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_154
timestamp -3599
transform 1 0 15272 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp -3599
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_169
timestamp -3599
transform 1 0 16652 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_175
timestamp -3599
transform 1 0 17204 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_180
timestamp 1636964856
transform 1 0 17664 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_192
timestamp 1636964856
transform 1 0 18768 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_204
timestamp 1636964856
transform 1 0 19872 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_216
timestamp -3599
transform 1 0 20976 0 -1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1636964856
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_237
timestamp 1636964856
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_249
timestamp 1636964856
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_261
timestamp -3599
transform 1 0 25116 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_265
timestamp -3599
transform 1 0 25484 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1636964856
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1636964856
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp -3599
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_29
timestamp -3599
transform 1 0 3772 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_37
timestamp -3599
transform 1 0 4508 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_43
timestamp -3599
transform 1 0 5060 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_48
timestamp -3599
transform 1 0 5520 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_57
timestamp -3599
transform 1 0 6348 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_66
timestamp -3599
transform 1 0 7176 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_74
timestamp -3599
transform 1 0 7912 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp -3599
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_85
timestamp -3599
transform 1 0 8924 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_93
timestamp -3599
transform 1 0 9660 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_100
timestamp -3599
transform 1 0 10304 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_105
timestamp -3599
transform 1 0 10764 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_112
timestamp -3599
transform 1 0 11408 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_121
timestamp -3599
transform 1 0 12236 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_128
timestamp -3599
transform 1 0 12880 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_135
timestamp -3599
transform 1 0 13524 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp -3599
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_141
timestamp -3599
transform 1 0 14076 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_146
timestamp -3599
transform 1 0 14536 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_155
timestamp -3599
transform 1 0 15364 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_159
timestamp -3599
transform 1 0 15732 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_168
timestamp -3599
transform 1 0 16560 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_175
timestamp -3599
transform 1 0 17204 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_182
timestamp -3599
transform 1 0 17848 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_189
timestamp -3599
transform 1 0 18492 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp -3599
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1636964856
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_209
timestamp 1636964856
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_221
timestamp 1636964856
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_233
timestamp 1636964856
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp -3599
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp -3599
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1636964856
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_265
timestamp -3599
transform 1 0 25484 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1636964856
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_15
timestamp -3599
transform 1 0 2484 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_28
timestamp -3599
transform 1 0 3680 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_37
timestamp -3599
transform 1 0 4508 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_44
timestamp -3599
transform 1 0 5152 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_53
timestamp -3599
transform 1 0 5980 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_29_57
timestamp -3599
transform 1 0 6348 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_61
timestamp -3599
transform 1 0 6716 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_70
timestamp -3599
transform 1 0 7544 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_77
timestamp -3599
transform 1 0 8188 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_82
timestamp -3599
transform 1 0 8648 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_91
timestamp -3599
transform 1 0 9476 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_100
timestamp -3599
transform 1 0 10304 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_106
timestamp -3599
transform 1 0 10856 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp -3599
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_113
timestamp -3599
transform 1 0 11500 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_122
timestamp -3599
transform 1 0 12328 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_130
timestamp -3599
transform 1 0 13064 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_136
timestamp -3599
transform 1 0 13616 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_147
timestamp 1636964856
transform 1 0 14628 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_159
timestamp -3599
transform 1 0 15732 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp -3599
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_169
timestamp -3599
transform 1 0 16652 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_173
timestamp -3599
transform 1 0 17020 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_194
timestamp -3599
transform 1 0 18952 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_214
timestamp -3599
transform 1 0 20792 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_222
timestamp -3599
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1636964856
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_237
timestamp 1636964856
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_249
timestamp 1636964856
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_261
timestamp -3599
transform 1 0 25116 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_265
timestamp -3599
transform 1 0 25484 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1636964856
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1636964856
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp -3599
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_29
timestamp -3599
transform 1 0 3772 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_37
timestamp -3599
transform 1 0 4508 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_42
timestamp -3599
transform 1 0 4968 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_47
timestamp -3599
transform 1 0 5428 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_55
timestamp -3599
transform 1 0 6164 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_64
timestamp -3599
transform 1 0 6992 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_71
timestamp -3599
transform 1 0 7636 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_78
timestamp -3599
transform 1 0 8280 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp -3599
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_85
timestamp -3599
transform 1 0 8924 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_92
timestamp -3599
transform 1 0 9568 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_99
timestamp -3599
transform 1 0 10212 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_104
timestamp -3599
transform 1 0 10672 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_109
timestamp -3599
transform 1 0 11132 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_116
timestamp -3599
transform 1 0 11776 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_125
timestamp -3599
transform 1 0 12604 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_132
timestamp -3599
transform 1 0 13248 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp -3599
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_141
timestamp -3599
transform 1 0 14076 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_151
timestamp -3599
transform 1 0 14996 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_30_158
timestamp -3599
transform 1 0 15640 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_167
timestamp -3599
transform 1 0 16468 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_174
timestamp -3599
transform 1 0 17112 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_186
timestamp -3599
transform 1 0 18216 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_191
timestamp -3599
transform 1 0 18676 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp -3599
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1636964856
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_209
timestamp 1636964856
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_221
timestamp 1636964856
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_233
timestamp 1636964856
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp -3599
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp -3599
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_253
timestamp 1636964856
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_265
timestamp -3599
transform 1 0 25484 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1636964856
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_15
timestamp -3599
transform 1 0 2484 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_24
timestamp -3599
transform 1 0 3312 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_33
timestamp -3599
transform 1 0 4140 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_41
timestamp -3599
transform 1 0 4876 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_48
timestamp -3599
transform 1 0 5520 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_53
timestamp -3599
transform 1 0 5980 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_31_57
timestamp -3599
transform 1 0 6348 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_67
timestamp -3599
transform 1 0 7268 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_71
timestamp 1636964856
transform 1 0 7636 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_83
timestamp -3599
transform 1 0 8740 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_88
timestamp -3599
transform 1 0 9200 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_95
timestamp -3599
transform 1 0 9844 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_104
timestamp -3599
transform 1 0 10672 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp -3599
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_113
timestamp -3599
transform 1 0 11500 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_122
timestamp -3599
transform 1 0 12328 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_128
timestamp -3599
transform 1 0 12880 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_138
timestamp -3599
transform 1 0 13800 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_143
timestamp -3599
transform 1 0 14260 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_151
timestamp -3599
transform 1 0 14996 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_159
timestamp -3599
transform 1 0 15732 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp -3599
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_169
timestamp -3599
transform 1 0 16652 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_177
timestamp -3599
transform 1 0 17388 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_186
timestamp 1636964856
transform 1 0 18216 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_198
timestamp 1636964856
transform 1 0 19320 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_210
timestamp 1636964856
transform 1 0 20424 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_222
timestamp -3599
transform 1 0 21528 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_225
timestamp 1636964856
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_237
timestamp 1636964856
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_249
timestamp 1636964856
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_261
timestamp -3599
transform 1 0 25116 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_265
timestamp -3599
transform 1 0 25484 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1636964856
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_15
timestamp -3599
transform 1 0 2484 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_23
timestamp -3599
transform 1 0 3220 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp -3599
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_29
timestamp -3599
transform 1 0 3772 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_37
timestamp -3599
transform 1 0 4508 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_43
timestamp -3599
transform 1 0 5060 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_48
timestamp -3599
transform 1 0 5520 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_53
timestamp -3599
transform 1 0 5980 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_63
timestamp -3599
transform 1 0 6900 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_74
timestamp -3599
transform 1 0 7912 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_82
timestamp -3599
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_85
timestamp -3599
transform 1 0 8924 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_92
timestamp -3599
transform 1 0 9568 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_96
timestamp -3599
transform 1 0 9936 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_104
timestamp -3599
transform 1 0 10672 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_108
timestamp -3599
transform 1 0 11040 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_118
timestamp -3599
transform 1 0 11960 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_127
timestamp -3599
transform 1 0 12788 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_132
timestamp -3599
transform 1 0 13248 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_141
timestamp -3599
transform 1 0 14076 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_149
timestamp -3599
transform 1 0 14812 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_155
timestamp 1636964856
transform 1 0 15364 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_167
timestamp -3599
transform 1 0 16468 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_173
timestamp -3599
transform 1 0 17020 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_178
timestamp -3599
transform 1 0 17480 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_183
timestamp 1636964856
transform 1 0 17940 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp -3599
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1636964856
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_209
timestamp 1636964856
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_221
timestamp 1636964856
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_233
timestamp 1636964856
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp -3599
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp -3599
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1636964856
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_265
timestamp -3599
transform 1 0 25484 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1636964856
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1636964856
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_27
timestamp -3599
transform 1 0 3588 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_37
timestamp -3599
transform 1 0 4508 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_41
timestamp -3599
transform 1 0 4876 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_47
timestamp -3599
transform 1 0 5428 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_52
timestamp -3599
transform 1 0 5888 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_57
timestamp -3599
transform 1 0 6348 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_61
timestamp -3599
transform 1 0 6716 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_65
timestamp -3599
transform 1 0 7084 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_70
timestamp -3599
transform 1 0 7544 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_79
timestamp -3599
transform 1 0 8372 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_83
timestamp -3599
transform 1 0 8740 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_90
timestamp -3599
transform 1 0 9384 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_97
timestamp -3599
transform 1 0 10028 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp -3599
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_113
timestamp -3599
transform 1 0 11500 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_122
timestamp -3599
transform 1 0 12328 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_126
timestamp -3599
transform 1 0 12696 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_132
timestamp -3599
transform 1 0 13248 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_140
timestamp -3599
transform 1 0 13984 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_149
timestamp -3599
transform 1 0 14812 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_162
timestamp -3599
transform 1 0 16008 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp -3599
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_169
timestamp -3599
transform 1 0 16652 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_177
timestamp 1636964856
transform 1 0 17388 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_189
timestamp 1636964856
transform 1 0 18492 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_201
timestamp 1636964856
transform 1 0 19596 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_213
timestamp -3599
transform 1 0 20700 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_221
timestamp -3599
transform 1 0 21436 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1636964856
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_237
timestamp 1636964856
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_249
timestamp 1636964856
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_261
timestamp -3599
transform 1 0 25116 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_265
timestamp -3599
transform 1 0 25484 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1636964856
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1636964856
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp -3599
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_29
timestamp -3599
transform 1 0 3772 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_33
timestamp -3599
transform 1 0 4140 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_41
timestamp -3599
transform 1 0 4876 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_50
timestamp -3599
transform 1 0 5704 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_56
timestamp -3599
transform 1 0 6256 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_60
timestamp -3599
transform 1 0 6624 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_64
timestamp -3599
transform 1 0 6992 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_73
timestamp -3599
transform 1 0 7820 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_82
timestamp -3599
transform 1 0 8648 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_85
timestamp -3599
transform 1 0 8924 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_91
timestamp -3599
transform 1 0 9476 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_98
timestamp -3599
transform 1 0 10120 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_103
timestamp -3599
transform 1 0 10580 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_34_116
timestamp -3599
transform 1 0 11776 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_121
timestamp -3599
transform 1 0 12236 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_130
timestamp -3599
transform 1 0 13064 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp -3599
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_141
timestamp -3599
transform 1 0 14076 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_145
timestamp -3599
transform 1 0 14444 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_154
timestamp -3599
transform 1 0 15272 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_161
timestamp -3599
transform 1 0 15916 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_168
timestamp -3599
transform 1 0 16560 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_173
timestamp -3599
transform 1 0 17020 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_178
timestamp 1636964856
transform 1 0 17480 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_190
timestamp -3599
transform 1 0 18584 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1636964856
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_209
timestamp 1636964856
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_221
timestamp 1636964856
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_233
timestamp 1636964856
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp -3599
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp -3599
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1636964856
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_265
timestamp -3599
transform 1 0 25484 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1636964856
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1636964856
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_27
timestamp -3599
transform 1 0 3588 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_29
timestamp -3599
transform 1 0 3772 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_35
timestamp -3599
transform 1 0 4324 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_42
timestamp -3599
transform 1 0 4968 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_49
timestamp -3599
transform 1 0 5612 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_54
timestamp -3599
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_57
timestamp -3599
transform 1 0 6348 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_61
timestamp -3599
transform 1 0 6716 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_67
timestamp -3599
transform 1 0 7268 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_75
timestamp -3599
transform 1 0 8004 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_35_83
timestamp -3599
transform 1 0 8740 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_85
timestamp -3599
transform 1 0 8924 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_90
timestamp -3599
transform 1 0 9384 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_95
timestamp -3599
transform 1 0 9844 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_100
timestamp 1636964856
transform 1 0 10304 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_113
timestamp -3599
transform 1 0 11500 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_120
timestamp -3599
transform 1 0 12144 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_127
timestamp 1636964856
transform 1 0 12788 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_139
timestamp -3599
transform 1 0 13892 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_141
timestamp -3599
transform 1 0 14076 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_147
timestamp -3599
transform 1 0 14628 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_152
timestamp -3599
transform 1 0 15088 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_157
timestamp -3599
transform 1 0 15548 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_164
timestamp -3599
transform 1 0 16192 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1636964856
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1636964856
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_193
timestamp -3599
transform 1 0 18860 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_197
timestamp 1636964856
transform 1 0 19228 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_209
timestamp 1636964856
transform 1 0 20332 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_221
timestamp -3599
transform 1 0 21436 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_225
timestamp 1636964856
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_237
timestamp 1636964856
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_249
timestamp -3599
transform 1 0 24012 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_253
timestamp 1636964856
transform 1 0 24380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_265
timestamp -3599
transform 1 0 25484 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_36
timestamp -3599
transform 1 0 1104 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp -3599
transform -1 0 25852 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_37
timestamp -3599
transform 1 0 1104 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp -3599
transform -1 0 25852 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_38
timestamp -3599
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp -3599
transform -1 0 25852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_39
timestamp -3599
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp -3599
transform -1 0 25852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_40
timestamp -3599
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp -3599
transform -1 0 25852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_41
timestamp -3599
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp -3599
transform -1 0 25852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_42
timestamp -3599
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp -3599
transform -1 0 25852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_43
timestamp -3599
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp -3599
transform -1 0 25852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_44
timestamp -3599
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp -3599
transform -1 0 25852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_45
timestamp -3599
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp -3599
transform -1 0 25852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_46
timestamp -3599
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp -3599
transform -1 0 25852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_47
timestamp -3599
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp -3599
transform -1 0 25852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_48
timestamp -3599
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp -3599
transform -1 0 25852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_49
timestamp -3599
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp -3599
transform -1 0 25852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_50
timestamp -3599
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp -3599
transform -1 0 25852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_51
timestamp -3599
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp -3599
transform -1 0 25852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_52
timestamp -3599
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp -3599
transform -1 0 25852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_53
timestamp -3599
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp -3599
transform -1 0 25852 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_54
timestamp -3599
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp -3599
transform -1 0 25852 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_55
timestamp -3599
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp -3599
transform -1 0 25852 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_56
timestamp -3599
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp -3599
transform -1 0 25852 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_57
timestamp -3599
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp -3599
transform -1 0 25852 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_58
timestamp -3599
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp -3599
transform -1 0 25852 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_59
timestamp -3599
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp -3599
transform -1 0 25852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_60
timestamp -3599
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp -3599
transform -1 0 25852 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_61
timestamp -3599
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp -3599
transform -1 0 25852 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_62
timestamp -3599
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp -3599
transform -1 0 25852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_63
timestamp -3599
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp -3599
transform -1 0 25852 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_64
timestamp -3599
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp -3599
transform -1 0 25852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_65
timestamp -3599
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp -3599
transform -1 0 25852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_66
timestamp -3599
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp -3599
transform -1 0 25852 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_67
timestamp -3599
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp -3599
transform -1 0 25852 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_68
timestamp -3599
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp -3599
transform -1 0 25852 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_69
timestamp -3599
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp -3599
transform -1 0 25852 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_70
timestamp -3599
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp -3599
transform -1 0 25852 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_71
timestamp -3599
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp -3599
transform -1 0 25852 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[0\].id.delaybuf0
timestamp -3599
transform 1 0 15364 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[0\].id.delaybuf1
timestamp -3599
transform -1 0 9384 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[0\].id.delayen0
timestamp -3599
transform 1 0 8004 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[0\].id.delayen1
timestamp -3599
transform 1 0 9016 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[0\].id.delayenb0
timestamp -3599
transform 1 0 7176 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_1  ringosc.dstage\[0\].id.delayenb1
timestamp -3599
transform 1 0 9568 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  ringosc.dstage\[0\].id.delayint0
timestamp -3599
transform -1 0 9844 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[1\].id.delaybuf0
timestamp -3599
transform -1 0 6992 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[1\].id.delaybuf1
timestamp -3599
transform 1 0 10304 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[1\].id.delayen0
timestamp -3599
transform -1 0 8372 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[1\].id.delayen1
timestamp -3599
transform 1 0 8280 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[1\].id.delayenb0
timestamp -3599
transform -1 0 8004 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_1  ringosc.dstage\[1\].id.delayenb1
timestamp -3599
transform -1 0 10120 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  ringosc.dstage\[1\].id.delayint0
timestamp -3599
transform -1 0 10304 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[2\].id.delaybuf0
timestamp -3599
transform 1 0 7268 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[2\].id.delaybuf1
timestamp -3599
transform 1 0 8464 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[2\].id.delayen0
timestamp -3599
transform -1 0 7544 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[2\].id.delayen1
timestamp -3599
transform 1 0 7176 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[2\].id.delayenb0
timestamp -3599
transform 1 0 6532 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_1  ringosc.dstage\[2\].id.delayenb1
timestamp -3599
transform -1 0 8280 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  ringosc.dstage\[2\].id.delayint0
timestamp -3599
transform 1 0 6440 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[3\].id.delaybuf0
timestamp -3599
transform 1 0 6716 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[3\].id.delaybuf1
timestamp -3599
transform 1 0 7084 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[3\].id.delayen0
timestamp -3599
transform 1 0 5704 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[3\].id.delayen1
timestamp -3599
transform 1 0 6440 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[3\].id.delayenb0
timestamp -3599
transform 1 0 5336 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_1  ringosc.dstage\[3\].id.delayenb1
timestamp -3599
transform 1 0 5704 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  ringosc.dstage\[3\].id.delayint0
timestamp -3599
transform -1 0 6624 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[4\].id.delaybuf0
timestamp -3599
transform 1 0 5244 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[4\].id.delaybuf1
timestamp -3599
transform 1 0 4784 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[4\].id.delayen0
timestamp -3599
transform 1 0 3864 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[4\].id.delayen1
timestamp -3599
transform -1 0 5152 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[4\].id.delayenb0
timestamp -3599
transform 1 0 3036 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_1  ringosc.dstage\[4\].id.delayenb1
timestamp -3599
transform -1 0 4508 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  ringosc.dstage\[4\].id.delayint0
timestamp -3599
transform -1 0 4968 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[5\].id.delaybuf0
timestamp -3599
transform -1 0 5428 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[5\].id.delaybuf1
timestamp -3599
transform 1 0 5704 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[5\].id.delayen0
timestamp -3599
transform -1 0 4508 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[5\].id.delayen1
timestamp -3599
transform 1 0 5060 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[5\].id.delayenb0
timestamp -3599
transform 1 0 3496 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_1  ringosc.dstage\[5\].id.delayenb1
timestamp -3599
transform 1 0 2852 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  ringosc.dstage\[5\].id.delayint0
timestamp -3599
transform 1 0 3312 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[6\].id.delaybuf0
timestamp -3599
transform -1 0 5520 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[6\].id.delaybuf1
timestamp -3599
transform 1 0 5796 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[6\].id.delayen0
timestamp -3599
transform 1 0 5060 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[6\].id.delayen1
timestamp -3599
transform 1 0 4968 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[6\].id.delayenb0
timestamp -3599
transform 1 0 4232 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_1  ringosc.dstage\[6\].id.delayenb1
timestamp -3599
transform 1 0 5152 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  ringosc.dstage\[6\].id.delayint0
timestamp -3599
transform -1 0 6716 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[7\].id.delaybuf0
timestamp -3599
transform -1 0 6256 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[7\].id.delaybuf1
timestamp -3599
transform -1 0 12236 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[7\].id.delayen0
timestamp -3599
transform 1 0 13248 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[7\].id.delayen1
timestamp -3599
transform 1 0 11684 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[7\].id.delayenb0
timestamp -3599
transform -1 0 13064 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_1  ringosc.dstage\[7\].id.delayenb1
timestamp -3599
transform 1 0 12328 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  ringosc.dstage\[7\].id.delayint0
timestamp -3599
transform 1 0 12972 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[8\].id.delaybuf0
timestamp -3599
transform -1 0 15088 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[8\].id.delaybuf1
timestamp -3599
transform 1 0 14168 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[8\].id.delayen0
timestamp -3599
transform 1 0 14628 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[8\].id.delayen1
timestamp -3599
transform -1 0 14628 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[8\].id.delayenb0
timestamp -3599
transform 1 0 14168 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_1  ringosc.dstage\[8\].id.delayenb1
timestamp -3599
transform -1 0 15916 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  ringosc.dstage\[8\].id.delayint0
timestamp -3599
transform -1 0 15548 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[9\].id.delaybuf0
timestamp -3599
transform -1 0 16468 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[9\].id.delaybuf1
timestamp -3599
transform 1 0 17204 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[9\].id.delayen0
timestamp -3599
transform -1 0 17388 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[9\].id.delayen1
timestamp -3599
transform 1 0 15732 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[9\].id.delayenb0
timestamp -3599
transform 1 0 15364 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_1  ringosc.dstage\[9\].id.delayenb1
timestamp -3599
transform 1 0 16100 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  ringosc.dstage\[9\].id.delayint0
timestamp -3599
transform -1 0 17020 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[10\].id.delaybuf0
timestamp -3599
transform -1 0 17020 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[10\].id.delaybuf1
timestamp -3599
transform 1 0 17204 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[10\].id.delayen0
timestamp -3599
transform 1 0 17572 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[10\].id.delayen1
timestamp -3599
transform 1 0 16652 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[10\].id.delayenb0
timestamp -3599
transform 1 0 16744 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_1  ringosc.dstage\[10\].id.delayenb1
timestamp -3599
transform 1 0 16008 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  ringosc.dstage\[10\].id.delayint0
timestamp -3599
transform 1 0 17664 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[11\].id.delaybuf0
timestamp -3599
transform 1 0 17848 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[11\].id.delaybuf1
timestamp -3599
transform 1 0 18400 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_8  ringosc.dstage\[11\].id.delayen0
timestamp -3599
transform -1 0 20792 0 -1 17408
box -38 -48 1694 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[11\].id.delayen1
timestamp -3599
transform 1 0 18032 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[11\].id.delayenb0
timestamp -3599
transform 1 0 17296 0 -1 17408
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_1  ringosc.dstage\[11\].id.delayenb1
timestamp -3599
transform 1 0 17388 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[11\].id.delayint0
timestamp -3599
transform 1 0 18676 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  ringosc.ibufp00
timestamp -3599
transform 1 0 16652 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_8  ringosc.ibufp01
timestamp -3599
transform 1 0 16744 0 -1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__clkinv_2  ringosc.ibufp10
timestamp -3599
transform -1 0 5060 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_4  ringosc.ibufp11
timestamp -3599
transform -1 0 4508 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__conb_1  ringosc.iss.const1
timestamp -3599
transform -1 0 16376 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  ringosc.iss.ctrlen0
timestamp -3599
transform 1 0 14812 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.iss.delaybuf0
timestamp -3599
transform 1 0 17388 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_4  ringosc.iss.delayen0
timestamp -3599
transform 1 0 15548 0 1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__einvp_1  ringosc.iss.delayen1
timestamp -3599
transform 1 0 16744 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_4  ringosc.iss.delayenb0
timestamp -3599
transform 1 0 15456 0 -1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__einvn_1  ringosc.iss.delayenb1
timestamp -3599
transform 1 0 16744 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  ringosc.iss.delayint0
timestamp -3599
transform -1 0 17020 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_4  ringosc.iss.reseten0
timestamp -3599
transform 1 0 15456 0 -1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_72
timestamp -3599
transform 1 0 3680 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_73
timestamp -3599
transform 1 0 6256 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_74
timestamp -3599
transform 1 0 8832 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_75
timestamp -3599
transform 1 0 11408 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_76
timestamp -3599
transform 1 0 13984 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_77
timestamp -3599
transform 1 0 16560 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_78
timestamp -3599
transform 1 0 19136 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_79
timestamp -3599
transform 1 0 21712 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_80
timestamp -3599
transform 1 0 24288 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_81
timestamp -3599
transform 1 0 6256 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_82
timestamp -3599
transform 1 0 11408 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_83
timestamp -3599
transform 1 0 16560 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_84
timestamp -3599
transform 1 0 21712 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_85
timestamp -3599
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_86
timestamp -3599
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_87
timestamp -3599
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_88
timestamp -3599
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_89
timestamp -3599
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_90
timestamp -3599
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_91
timestamp -3599
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_92
timestamp -3599
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_93
timestamp -3599
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_94
timestamp -3599
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_95
timestamp -3599
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_96
timestamp -3599
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_97
timestamp -3599
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_98
timestamp -3599
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_99
timestamp -3599
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_100
timestamp -3599
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_101
timestamp -3599
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_102
timestamp -3599
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_103
timestamp -3599
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_104
timestamp -3599
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_105
timestamp -3599
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_106
timestamp -3599
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_107
timestamp -3599
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_108
timestamp -3599
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_109
timestamp -3599
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_110
timestamp -3599
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_111
timestamp -3599
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_112
timestamp -3599
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_113
timestamp -3599
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_114
timestamp -3599
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_115
timestamp -3599
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_116
timestamp -3599
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_117
timestamp -3599
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_118
timestamp -3599
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_119
timestamp -3599
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_120
timestamp -3599
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_121
timestamp -3599
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_122
timestamp -3599
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_123
timestamp -3599
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_124
timestamp -3599
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_125
timestamp -3599
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_126
timestamp -3599
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_127
timestamp -3599
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_128
timestamp -3599
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_129
timestamp -3599
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_130
timestamp -3599
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_131
timestamp -3599
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_132
timestamp -3599
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_133
timestamp -3599
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_134
timestamp -3599
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_135
timestamp -3599
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_136
timestamp -3599
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_137
timestamp -3599
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_138
timestamp -3599
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_139
timestamp -3599
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_140
timestamp -3599
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_141
timestamp -3599
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_142
timestamp -3599
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_143
timestamp -3599
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_144
timestamp -3599
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_145
timestamp -3599
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_146
timestamp -3599
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_147
timestamp -3599
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_148
timestamp -3599
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_149
timestamp -3599
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_150
timestamp -3599
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_151
timestamp -3599
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_152
timestamp -3599
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_153
timestamp -3599
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_154
timestamp -3599
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_155
timestamp -3599
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_156
timestamp -3599
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_157
timestamp -3599
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_158
timestamp -3599
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_159
timestamp -3599
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_160
timestamp -3599
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_161
timestamp -3599
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_162
timestamp -3599
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_163
timestamp -3599
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_164
timestamp -3599
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_165
timestamp -3599
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_166
timestamp -3599
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_167
timestamp -3599
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_168
timestamp -3599
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_169
timestamp -3599
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_170
timestamp -3599
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_171
timestamp -3599
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_172
timestamp -3599
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_173
timestamp -3599
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_174
timestamp -3599
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_175
timestamp -3599
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_176
timestamp -3599
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_177
timestamp -3599
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_178
timestamp -3599
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_179
timestamp -3599
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_180
timestamp -3599
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_181
timestamp -3599
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_182
timestamp -3599
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_183
timestamp -3599
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_184
timestamp -3599
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_185
timestamp -3599
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_186
timestamp -3599
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_187
timestamp -3599
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_188
timestamp -3599
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_189
timestamp -3599
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_190
timestamp -3599
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_191
timestamp -3599
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_192
timestamp -3599
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_193
timestamp -3599
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_194
timestamp -3599
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_195
timestamp -3599
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_196
timestamp -3599
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_197
timestamp -3599
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_198
timestamp -3599
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_199
timestamp -3599
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_200
timestamp -3599
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_201
timestamp -3599
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_202
timestamp -3599
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_203
timestamp -3599
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_204
timestamp -3599
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_205
timestamp -3599
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_206
timestamp -3599
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_207
timestamp -3599
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_208
timestamp -3599
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_209
timestamp -3599
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_210
timestamp -3599
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_211
timestamp -3599
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_212
timestamp -3599
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_213
timestamp -3599
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_214
timestamp -3599
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_215
timestamp -3599
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_216
timestamp -3599
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_217
timestamp -3599
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_218
timestamp -3599
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_219
timestamp -3599
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_220
timestamp -3599
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_221
timestamp -3599
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_222
timestamp -3599
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_223
timestamp -3599
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_224
timestamp -3599
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_225
timestamp -3599
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_226
timestamp -3599
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_227
timestamp -3599
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_228
timestamp -3599
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_229
timestamp -3599
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_230
timestamp -3599
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_231
timestamp -3599
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_232
timestamp -3599
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_233
timestamp -3599
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_234
timestamp -3599
transform 1 0 3680 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_235
timestamp -3599
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_236
timestamp -3599
transform 1 0 8832 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_237
timestamp -3599
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_238
timestamp -3599
transform 1 0 13984 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_239
timestamp -3599
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_240
timestamp -3599
transform 1 0 19136 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_241
timestamp -3599
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_242
timestamp -3599
transform 1 0 24288 0 -1 20672
box -38 -48 130 592
<< labels >>
flabel metal4 s 8208 1040 8528 20720 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 16208 1040 16528 20720 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 24208 1040 24528 20720 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4208 1040 4528 20720 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 12208 1040 12528 20720 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 20208 1040 20528 20720 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 1096 800 1216 0 FreeSans 480 0 0 0 clockp[0]
port 2 nsew signal output
flabel metal3 s 0 2184 800 2304 0 FreeSans 480 0 0 0 clockp[1]
port 3 nsew signal output
flabel metal3 s 0 13064 800 13184 0 FreeSans 480 0 0 0 dco
port 4 nsew signal input
flabel metal3 s 0 3272 800 3392 0 FreeSans 480 0 0 0 div[0]
port 5 nsew signal input
flabel metal3 s 0 4360 800 4480 0 FreeSans 480 0 0 0 div[1]
port 6 nsew signal input
flabel metal3 s 0 5448 800 5568 0 FreeSans 480 0 0 0 div[2]
port 7 nsew signal input
flabel metal3 s 0 6536 800 6656 0 FreeSans 480 0 0 0 div[3]
port 8 nsew signal input
flabel metal3 s 0 7624 800 7744 0 FreeSans 480 0 0 0 div[4]
port 9 nsew signal input
flabel metal3 s 0 8712 800 8832 0 FreeSans 480 0 0 0 div[5]
port 10 nsew signal input
flabel metal3 s 0 9800 800 9920 0 FreeSans 480 0 0 0 div[6]
port 11 nsew signal input
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 div[7]
port 12 nsew signal input
flabel metal3 s 0 11976 800 12096 0 FreeSans 480 0 0 0 enable
port 13 nsew signal input
flabel metal3 s 0 14152 800 14272 0 FreeSans 480 0 0 0 ext_trim[0]
port 14 nsew signal input
flabel metal2 s 7378 21200 7434 22000 0 FreeSans 224 90 0 0 ext_trim[10]
port 15 nsew signal input
flabel metal2 s 9402 21200 9458 22000 0 FreeSans 224 90 0 0 ext_trim[11]
port 16 nsew signal input
flabel metal2 s 11426 21200 11482 22000 0 FreeSans 224 90 0 0 ext_trim[12]
port 17 nsew signal input
flabel metal2 s 13450 21200 13506 22000 0 FreeSans 224 90 0 0 ext_trim[13]
port 18 nsew signal input
flabel metal2 s 15474 21200 15530 22000 0 FreeSans 224 90 0 0 ext_trim[14]
port 19 nsew signal input
flabel metal2 s 17498 21200 17554 22000 0 FreeSans 224 90 0 0 ext_trim[15]
port 20 nsew signal input
flabel metal2 s 19522 21200 19578 22000 0 FreeSans 224 90 0 0 ext_trim[16]
port 21 nsew signal input
flabel metal2 s 21546 21200 21602 22000 0 FreeSans 224 90 0 0 ext_trim[17]
port 22 nsew signal input
flabel metal2 s 23570 21200 23626 22000 0 FreeSans 224 90 0 0 ext_trim[18]
port 23 nsew signal input
flabel metal2 s 25594 21200 25650 22000 0 FreeSans 224 90 0 0 ext_trim[19]
port 24 nsew signal input
flabel metal3 s 0 15240 800 15360 0 FreeSans 480 0 0 0 ext_trim[1]
port 25 nsew signal input
flabel metal3 s 26200 19592 27000 19712 0 FreeSans 480 0 0 0 ext_trim[20]
port 26 nsew signal input
flabel metal3 s 26200 16056 27000 16176 0 FreeSans 480 0 0 0 ext_trim[21]
port 27 nsew signal input
flabel metal3 s 26200 12520 27000 12640 0 FreeSans 480 0 0 0 ext_trim[22]
port 28 nsew signal input
flabel metal3 s 26200 8984 27000 9104 0 FreeSans 480 0 0 0 ext_trim[23]
port 29 nsew signal input
flabel metal3 s 26200 5448 27000 5568 0 FreeSans 480 0 0 0 ext_trim[24]
port 30 nsew signal input
flabel metal3 s 26200 1912 27000 2032 0 FreeSans 480 0 0 0 ext_trim[25]
port 31 nsew signal input
flabel metal3 s 0 16328 800 16448 0 FreeSans 480 0 0 0 ext_trim[2]
port 32 nsew signal input
flabel metal3 s 0 17416 800 17536 0 FreeSans 480 0 0 0 ext_trim[3]
port 33 nsew signal input
flabel metal3 s 0 18504 800 18624 0 FreeSans 480 0 0 0 ext_trim[4]
port 34 nsew signal input
flabel metal3 s 0 19592 800 19712 0 FreeSans 480 0 0 0 ext_trim[5]
port 35 nsew signal input
flabel metal3 s 0 20680 800 20800 0 FreeSans 480 0 0 0 ext_trim[6]
port 36 nsew signal input
flabel metal2 s 1306 21200 1362 22000 0 FreeSans 224 90 0 0 ext_trim[7]
port 37 nsew signal input
flabel metal2 s 3330 21200 3386 22000 0 FreeSans 224 90 0 0 ext_trim[8]
port 38 nsew signal input
flabel metal2 s 5354 21200 5410 22000 0 FreeSans 224 90 0 0 ext_trim[9]
port 39 nsew signal input
flabel metal2 s 20166 0 20222 800 0 FreeSans 224 90 0 0 osc
port 40 nsew signal input
flabel metal2 s 6734 0 6790 800 0 FreeSans 224 90 0 0 resetb
port 41 nsew signal input
rlabel metal1 13478 20672 13478 20672 0 VGND
rlabel metal1 13478 20128 13478 20128 0 VPWR
rlabel metal1 4508 15878 4508 15878 0 _000_
rlabel metal2 2990 15198 2990 15198 0 _001_
rlabel metal1 3220 15878 3220 15878 0 _002_
rlabel metal2 9798 11934 9798 11934 0 _003_
rlabel metal2 8142 15198 8142 15198 0 _004_
rlabel metal1 10166 13158 10166 13158 0 _005_
rlabel metal2 15502 13430 15502 13430 0 _006_
rlabel metal2 15042 13090 15042 13090 0 _007_
rlabel metal2 14950 11934 14950 11934 0 _008_
rlabel metal1 16613 11050 16613 11050 0 _009_
rlabel metal1 16889 12138 16889 12138 0 _010_
rlabel metal1 19274 12070 19274 12070 0 _011_
rlabel metal1 18439 11798 18439 11798 0 _012_
rlabel metal1 20700 8602 20700 8602 0 _013_
rlabel metal1 14536 4998 14536 4998 0 _014_
rlabel metal2 20470 2142 20470 2142 0 _015_
rlabel metal1 16422 2822 16422 2822 0 _016_
rlabel metal1 18216 6086 18216 6086 0 _017_
rlabel metal2 21022 4250 21022 4250 0 _018_
rlabel metal1 23039 7446 23039 7446 0 _019_
rlabel metal1 10718 8602 10718 8602 0 _020_
rlabel metal2 12650 10642 12650 10642 0 _021_
rlabel metal1 9667 10710 9667 10710 0 _022_
rlabel metal2 11086 10268 11086 10268 0 _023_
rlabel metal2 9338 10336 9338 10336 0 _024_
rlabel metal2 12006 9792 12006 9792 0 _025_
rlabel metal1 13425 7446 13425 7446 0 _026_
rlabel metal1 19918 4046 19918 4046 0 _027_
rlabel metal1 19097 3434 19097 3434 0 _028_
rlabel metal1 20654 5338 20654 5338 0 _029_
rlabel metal1 23644 3706 23644 3706 0 _030_
rlabel metal2 23690 6120 23690 6120 0 _031_
rlabel metal2 11178 3502 11178 3502 0 _032_
rlabel metal2 10626 3706 10626 3706 0 _033_
rlabel metal1 9200 4794 9200 4794 0 _034_
rlabel metal1 10120 6086 10120 6086 0 _035_
rlabel metal1 9023 8534 9023 8534 0 _036_
rlabel metal1 9706 6834 9706 6834 0 _037_
rlabel metal2 14398 2414 14398 2414 0 _038_
rlabel metal2 17526 2142 17526 2142 0 _039_
rlabel metal1 13885 2346 13885 2346 0 _040_
rlabel metal1 15916 7718 15916 7718 0 _041_
rlabel metal1 21903 6698 21903 6698 0 _042_
rlabel metal1 21942 8602 21942 8602 0 _043_
rlabel metal2 15502 9384 15502 9384 0 _044_
rlabel metal1 19274 10234 19274 10234 0 _045_
rlabel metal2 17710 9384 17710 9384 0 _046_
rlabel metal2 21206 10200 21206 10200 0 _047_
rlabel metal2 22770 10472 22770 10472 0 _048_
rlabel metal1 24472 9146 24472 9146 0 _049_
rlabel metal2 21114 3366 21114 3366 0 _050_
rlabel metal2 22034 3298 22034 3298 0 _051_
rlabel metal2 16514 3944 16514 3944 0 _052_
rlabel metal1 12611 2346 12611 2346 0 _053_
rlabel metal1 10679 2006 10679 2006 0 _054_
rlabel metal2 13018 4318 13018 4318 0 _055_
rlabel metal2 12650 5032 12650 5032 0 _056_
rlabel metal2 12006 6936 12006 6936 0 _057_
rlabel metal2 11914 8738 11914 8738 0 _058_
rlabel metal1 15226 8058 15226 8058 0 _059_
rlabel metal1 17894 6630 17894 6630 0 _060_
rlabel metal1 18499 7786 18499 7786 0 _061_
rlabel metal2 20378 7684 20378 7684 0 _062_
rlabel metal1 23177 4182 23177 4182 0 _063_
rlabel metal1 23506 8058 23506 8058 0 _064_
rlabel metal1 4600 3366 4600 3366 0 _065_
rlabel metal2 4186 2261 4186 2261 0 _066_
rlabel metal1 2898 3706 2898 3706 0 _067_
rlabel metal2 2806 5542 2806 5542 0 _068_
rlabel metal2 2806 6936 2806 6936 0 _069_
rlabel metal2 2806 8262 2806 8262 0 _070_
rlabel metal1 2576 10438 2576 10438 0 _071_
rlabel metal2 2622 11934 2622 11934 0 _072_
rlabel metal1 6394 11254 6394 11254 0 _073_
rlabel metal1 4186 15368 4186 15368 0 _074_
rlabel metal2 2714 14382 2714 14382 0 _075_
rlabel metal1 2070 14280 2070 14280 0 _076_
rlabel metal1 8464 12614 8464 12614 0 _077_
rlabel metal1 6992 14586 6992 14586 0 _078_
rlabel metal1 9936 13226 9936 13226 0 _079_
rlabel metal2 14398 14110 14398 14110 0 _080_
rlabel metal2 14490 13906 14490 13906 0 _081_
rlabel metal2 13386 11186 13386 11186 0 _082_
rlabel metal2 16974 11356 16974 11356 0 _083_
rlabel metal2 17250 12002 17250 12002 0 _084_
rlabel metal2 19550 11730 19550 11730 0 _085_
rlabel metal1 18032 11322 18032 11322 0 _086_
rlabel metal1 19780 8602 19780 8602 0 _087_
rlabel metal2 14398 4250 14398 4250 0 _088_
rlabel metal2 19090 2142 19090 2142 0 _089_
rlabel metal1 17710 2312 17710 2312 0 _090_
rlabel metal2 17250 5848 17250 5848 0 _091_
rlabel metal2 20746 4828 20746 4828 0 _092_
rlabel metal2 22678 7582 22678 7582 0 _093_
rlabel metal2 9614 9180 9614 9180 0 _094_
rlabel metal1 11858 11322 11858 11322 0 _095_
rlabel metal2 8142 10846 8142 10846 0 _096_
rlabel via1 9975 11322 9975 11322 0 _097_
rlabel metal2 7774 10370 7774 10370 0 _098_
rlabel metal1 10488 9690 10488 9690 0 _099_
rlabel metal1 13570 6970 13570 6970 0 _100_
rlabel metal1 18492 4182 18492 4182 0 _101_
rlabel metal2 17526 4012 17526 4012 0 _102_
rlabel metal2 19826 5916 19826 5916 0 _103_
rlabel metal2 23138 4930 23138 4930 0 _104_
rlabel metal1 23782 6222 23782 6222 0 _105_
rlabel metal2 9338 3230 9338 3230 0 _106_
rlabel metal1 9660 3434 9660 3434 0 _107_
rlabel metal2 9614 5678 9614 5678 0 _108_
rlabel metal1 9016 5610 9016 5610 0 _109_
rlabel metal2 7406 7684 7406 7684 0 _110_
rlabel metal2 8050 7582 8050 7582 0 _111_
rlabel metal1 14720 3366 14720 3366 0 _112_
rlabel metal2 17066 1700 17066 1700 0 _113_
rlabel metal1 15364 3026 15364 3026 0 _114_
rlabel metal2 15134 6052 15134 6052 0 _115_
rlabel metal2 21390 6630 21390 6630 0 _116_
rlabel metal2 22862 9180 22862 9180 0 _117_
rlabel metal2 14490 10030 14490 10030 0 _118_
rlabel metal2 18814 10132 18814 10132 0 _119_
rlabel metal1 17020 9622 17020 9622 0 _120_
rlabel metal1 20286 9962 20286 9962 0 _121_
rlabel metal2 22310 11016 22310 11016 0 _122_
rlabel metal1 23046 9486 23046 9486 0 _123_
rlabel metal1 11408 1530 11408 1530 0 _124_
rlabel metal1 11040 1530 11040 1530 0 _125_
rlabel metal1 12144 3706 12144 3706 0 _126_
rlabel metal2 11914 4964 11914 4964 0 _127_
rlabel metal1 11447 6970 11447 6970 0 _128_
rlabel metal2 12466 8704 12466 8704 0 _129_
rlabel metal2 15502 8670 15502 8670 0 _130_
rlabel metal2 18906 7582 18906 7582 0 _131_
rlabel metal2 16974 8092 16974 8092 0 _132_
rlabel metal1 21252 7922 21252 7922 0 _133_
rlabel metal2 23322 4794 23322 4794 0 _134_
rlabel metal1 23782 8058 23782 8058 0 _135_
rlabel metal1 5474 2006 5474 2006 0 _136_
rlabel metal2 3174 2142 3174 2142 0 _137_
rlabel metal1 2116 3706 2116 3706 0 _138_
rlabel metal1 1932 5270 1932 5270 0 _139_
rlabel metal1 1978 6426 1978 6426 0 _140_
rlabel metal2 1794 8670 1794 8670 0 _141_
rlabel metal1 1932 9690 1932 9690 0 _142_
rlabel metal1 2116 11322 2116 11322 0 _143_
rlabel metal2 5842 11934 5842 11934 0 _144_
rlabel via1 4001 11730 4001 11730 0 _145_
rlabel metal2 6578 9758 6578 9758 0 _146_
rlabel metal1 6578 9078 6578 9078 0 _147_
rlabel metal2 6762 9350 6762 9350 0 _148_
rlabel metal2 6486 10404 6486 10404 0 _149_
rlabel metal1 7130 9350 7130 9350 0 _150_
rlabel metal1 6440 10642 6440 10642 0 _151_
rlabel metal2 5566 8058 5566 8058 0 _152_
rlabel metal2 5750 7616 5750 7616 0 _153_
rlabel metal1 6164 7242 6164 7242 0 _154_
rlabel metal1 6210 7514 6210 7514 0 _155_
rlabel metal1 5980 7786 5980 7786 0 _156_
rlabel metal2 5290 5202 5290 5202 0 _157_
rlabel metal1 6440 5678 6440 5678 0 _158_
rlabel metal1 7268 5338 7268 5338 0 _159_
rlabel metal1 7728 4658 7728 4658 0 _160_
rlabel metal1 7774 5202 7774 5202 0 _161_
rlabel metal1 7038 5542 7038 5542 0 _162_
rlabel metal1 7498 1836 7498 1836 0 _163_
rlabel metal1 8832 1326 8832 1326 0 _164_
rlabel metal1 7452 2482 7452 2482 0 _165_
rlabel metal1 8096 1394 8096 1394 0 _166_
rlabel via1 7406 1394 7406 1394 0 _167_
rlabel metal2 8418 1700 8418 1700 0 _168_
rlabel metal2 7774 2788 7774 2788 0 _169_
rlabel metal2 7498 4284 7498 4284 0 _170_
rlabel metal1 8188 4114 8188 4114 0 _171_
rlabel metal1 8556 2618 8556 2618 0 _172_
rlabel metal1 7866 3570 7866 3570 0 _173_
rlabel metal2 7590 3706 7590 3706 0 _174_
rlabel metal1 7084 5134 7084 5134 0 _175_
rlabel metal1 6716 5066 6716 5066 0 _176_
rlabel metal1 6486 6290 6486 6290 0 _177_
rlabel metal1 5290 6256 5290 6256 0 _178_
rlabel metal2 5198 6562 5198 6562 0 _179_
rlabel metal1 5244 6630 5244 6630 0 _180_
rlabel metal1 6118 6256 6118 6256 0 _181_
rlabel metal1 5934 6324 5934 6324 0 _182_
rlabel metal1 5428 6154 5428 6154 0 _183_
rlabel metal2 6394 7140 6394 7140 0 _184_
rlabel metal1 5566 7956 5566 7956 0 _185_
rlabel metal1 6532 10438 6532 10438 0 _186_
rlabel metal1 5842 10506 5842 10506 0 _187_
rlabel metal2 4738 11271 4738 11271 0 _188_
rlabel metal1 5014 12172 5014 12172 0 _189_
rlabel metal2 4830 11798 4830 11798 0 _190_
rlabel metal2 5566 11628 5566 11628 0 _191_
rlabel metal1 16882 6290 16882 6290 0 _192_
rlabel metal1 14214 10506 14214 10506 0 _193_
rlabel metal1 4048 5134 4048 5134 0 _194_
rlabel metal2 6026 11764 6026 11764 0 _195_
rlabel metal1 4462 10642 4462 10642 0 _196_
rlabel metal1 3588 10778 3588 10778 0 _197_
rlabel metal1 2806 11186 2806 11186 0 _198_
rlabel metal1 3680 9622 3680 9622 0 _199_
rlabel metal1 2438 9554 2438 9554 0 _200_
rlabel viali 4816 7378 4816 7378 0 _201_
rlabel metal2 4462 7616 4462 7616 0 _202_
rlabel metal1 2438 8058 2438 8058 0 _203_
rlabel metal1 3818 6154 3818 6154 0 _204_
rlabel metal1 2806 6358 2806 6358 0 _205_
rlabel metal1 6854 5236 6854 5236 0 _206_
rlabel metal1 5244 5338 5244 5338 0 _207_
rlabel metal1 2254 5644 2254 5644 0 _208_
rlabel metal1 6486 3570 6486 3570 0 _209_
rlabel metal2 6670 3876 6670 3876 0 _210_
rlabel metal1 25070 7956 25070 7956 0 _211_
rlabel metal1 2438 3536 2438 3536 0 _212_
rlabel metal1 6578 1870 6578 1870 0 _213_
rlabel metal2 6854 1904 6854 1904 0 _214_
rlabel metal1 3542 2346 3542 2346 0 _215_
rlabel metal1 7590 5848 7590 5848 0 _216_
rlabel metal1 17204 4046 17204 4046 0 _217_
rlabel metal1 7912 1734 7912 1734 0 _218_
rlabel metal1 6992 1938 6992 1938 0 _219_
rlabel metal1 24288 7854 24288 7854 0 _220_
rlabel metal2 23414 5236 23414 5236 0 _221_
rlabel metal1 20792 7514 20792 7514 0 _222_
rlabel metal1 17204 8466 17204 8466 0 _223_
rlabel metal1 19504 7854 19504 7854 0 _224_
rlabel metal1 13202 6222 13202 6222 0 _225_
rlabel metal1 16146 8976 16146 8976 0 _226_
rlabel metal1 12742 8534 12742 8534 0 _227_
rlabel metal1 11868 6426 11868 6426 0 _228_
rlabel metal2 12098 5066 12098 5066 0 _229_
rlabel metal1 12604 3502 12604 3502 0 _230_
rlabel metal1 11454 2822 11454 2822 0 _231_
rlabel metal2 11822 1530 11822 1530 0 _232_
rlabel metal1 23598 10132 23598 10132 0 _233_
rlabel metal1 22678 9554 22678 9554 0 _234_
rlabel metal1 21988 11118 21988 11118 0 _235_
rlabel metal1 20332 11118 20332 11118 0 _236_
rlabel metal1 16882 10234 16882 10234 0 _237_
rlabel metal2 18998 9724 18998 9724 0 _238_
rlabel metal2 14950 10438 14950 10438 0 _239_
rlabel metal1 22770 9146 22770 9146 0 _240_
rlabel metal1 22632 6222 22632 6222 0 _241_
rlabel metal1 21758 6290 21758 6290 0 _242_
rlabel metal1 15456 5678 15456 5678 0 _243_
rlabel metal1 13754 3060 13754 3060 0 _244_
rlabel metal1 17434 1326 17434 1326 0 _245_
rlabel metal1 14398 3502 14398 3502 0 _246_
rlabel metal2 10350 5712 10350 5712 0 _247_
rlabel metal1 8326 6698 8326 6698 0 _248_
rlabel metal2 7774 7242 7774 7242 0 _249_
rlabel metal1 7866 6800 7866 6800 0 _250_
rlabel metal2 8234 5882 8234 5882 0 _251_
rlabel metal1 8602 10132 8602 10132 0 _252_
rlabel metal1 9660 4114 9660 4114 0 _253_
rlabel metal1 10166 5236 10166 5236 0 _254_
rlabel metal1 10074 5338 10074 5338 0 _255_
rlabel metal1 9890 4046 9890 4046 0 _256_
rlabel metal1 24564 6970 24564 6970 0 _257_
rlabel metal1 23736 4590 23736 4590 0 _258_
rlabel metal1 20240 6290 20240 6290 0 _259_
rlabel metal1 17802 4250 17802 4250 0 _260_
rlabel metal1 19044 4590 19044 4590 0 _261_
rlabel metal1 14168 6630 14168 6630 0 _262_
rlabel metal2 10442 9078 10442 9078 0 _263_
rlabel metal2 7958 10676 7958 10676 0 _264_
rlabel metal1 10396 10778 10396 10778 0 _265_
rlabel metal2 9062 10676 9062 10676 0 _266_
rlabel metal1 11592 10778 11592 10778 0 _267_
rlabel metal2 10718 8806 10718 8806 0 _268_
rlabel metal1 23184 6970 23184 6970 0 _269_
rlabel metal1 21666 5202 21666 5202 0 _270_
rlabel metal1 18906 5134 18906 5134 0 _271_
rlabel metal1 17802 5338 17802 5338 0 _272_
rlabel metal1 18078 2822 18078 2822 0 _273_
rlabel metal1 19090 2414 19090 2414 0 _274_
rlabel metal2 14214 4590 14214 4590 0 _275_
rlabel metal2 19550 8636 19550 8636 0 _276_
rlabel metal1 18032 11118 18032 11118 0 _277_
rlabel metal1 19596 11118 19596 11118 0 _278_
rlabel metal1 17434 11696 17434 11696 0 _279_
rlabel metal2 16790 11254 16790 11254 0 _280_
rlabel metal1 13432 10642 13432 10642 0 _281_
rlabel metal2 3634 8772 3634 8772 0 _282_
rlabel metal1 5290 8432 5290 8432 0 _283_
rlabel metal2 4646 9231 4646 9231 0 _284_
rlabel metal1 4048 9078 4048 9078 0 _285_
rlabel metal1 5566 9554 5566 9554 0 _286_
rlabel metal2 6118 9792 6118 9792 0 _287_
rlabel metal1 6808 9894 6808 9894 0 _288_
rlabel metal1 6716 10030 6716 10030 0 _289_
rlabel metal1 4784 9418 4784 9418 0 _290_
rlabel metal2 5382 9724 5382 9724 0 _291_
rlabel metal1 4830 9554 4830 9554 0 _292_
rlabel metal1 4232 8466 4232 8466 0 _293_
rlabel metal1 4784 8330 4784 8330 0 _294_
rlabel metal2 4738 7106 4738 7106 0 _295_
rlabel metal1 4531 4794 4531 4794 0 _296_
rlabel metal1 2346 4556 2346 4556 0 _297_
rlabel metal1 2530 4760 2530 4760 0 _298_
rlabel metal1 2661 4522 2661 4522 0 _299_
rlabel metal1 4324 5270 4324 5270 0 _300_
rlabel metal1 4600 3094 4600 3094 0 _301_
rlabel metal1 4922 1530 4922 1530 0 _302_
rlabel metal2 4922 2417 4922 2417 0 _303_
rlabel metal1 4324 3162 4324 3162 0 _304_
rlabel metal1 4462 4250 4462 4250 0 _305_
rlabel metal1 5152 5066 5152 5066 0 _306_
rlabel metal1 3956 12818 3956 12818 0 _307_
rlabel metal1 10994 14416 10994 14416 0 _308_
rlabel metal1 11040 13906 11040 13906 0 _309_
rlabel metal1 8464 13498 8464 13498 0 _310_
rlabel metal1 5934 12886 5934 12886 0 _311_
rlabel metal2 2162 14178 2162 14178 0 _312_
rlabel metal2 3542 14382 3542 14382 0 _313_
rlabel metal1 2438 13838 2438 13838 0 _314_
rlabel metal1 4554 13430 4554 13430 0 _315_
rlabel metal1 4554 12852 4554 12852 0 _316_
rlabel metal1 5750 12716 5750 12716 0 _317_
rlabel metal1 5842 13328 5842 13328 0 _318_
rlabel metal1 6808 13362 6808 13362 0 _319_
rlabel metal1 7590 14348 7590 14348 0 _320_
rlabel metal1 10350 13974 10350 13974 0 _321_
rlabel metal2 11270 13260 11270 13260 0 _322_
rlabel metal2 12926 14144 12926 14144 0 _323_
rlabel metal1 5394 2958 5394 2958 0 _324_
rlabel metal1 5244 3162 5244 3162 0 _325_
rlabel metal2 6394 12857 6394 12857 0 _326_
rlabel metal1 9706 14484 9706 14484 0 _327_
rlabel metal1 12006 16490 12006 16490 0 _328_
rlabel viali 8417 13906 8417 13906 0 _329_
rlabel metal1 6992 13294 6992 13294 0 _330_
rlabel metal1 8694 16626 8694 16626 0 _331_
rlabel metal2 13018 17748 13018 17748 0 _332_
rlabel via2 12650 18717 12650 18717 0 _333_
rlabel metal1 8188 16966 8188 16966 0 _334_
rlabel metal2 5750 14348 5750 14348 0 _335_
rlabel metal2 6486 13498 6486 13498 0 _336_
rlabel metal2 9522 13294 9522 13294 0 _337_
rlabel metal2 12834 13872 12834 13872 0 _338_
rlabel metal2 12006 14042 12006 14042 0 _339_
rlabel metal2 13386 13498 13386 13498 0 _340_
rlabel metal1 13984 13498 13984 13498 0 _341_
rlabel metal1 11408 12954 11408 12954 0 _342_
rlabel metal2 10534 13328 10534 13328 0 _343_
rlabel metal1 9706 12954 9706 12954 0 _344_
rlabel metal1 7682 13328 7682 13328 0 _345_
rlabel metal1 7452 13498 7452 13498 0 _346_
rlabel metal1 6900 14042 6900 14042 0 _347_
rlabel metal1 6210 12750 6210 12750 0 _348_
rlabel metal1 6808 12954 6808 12954 0 _349_
rlabel metal1 8004 12818 8004 12818 0 _350_
rlabel metal2 4002 14348 4002 14348 0 _351_
rlabel metal1 3220 13294 3220 13294 0 _352_
rlabel metal1 4462 14416 4462 14416 0 _353_
rlabel metal1 3634 14042 3634 14042 0 _354_
rlabel metal2 7130 19142 7130 19142 0 _355_
rlabel metal1 12558 18190 12558 18190 0 _356_
rlabel metal1 10810 16558 10810 16558 0 _357_
rlabel metal1 11684 16558 11684 16558 0 _358_
rlabel metal1 13386 16184 13386 16184 0 _359_
rlabel metal1 12466 18394 12466 18394 0 _360_
rlabel metal1 13754 18666 13754 18666 0 _361_
rlabel metal1 6256 18734 6256 18734 0 _362_
rlabel metal1 10258 18292 10258 18292 0 _363_
rlabel metal1 12558 16660 12558 16660 0 _364_
rlabel via2 11638 16779 11638 16779 0 _365_
rlabel metal2 11546 17306 11546 17306 0 _366_
rlabel metal2 12190 17408 12190 17408 0 _367_
rlabel metal1 8832 18734 8832 18734 0 _368_
rlabel metal1 8234 16218 8234 16218 0 _369_
rlabel metal2 10074 15538 10074 15538 0 _370_
rlabel viali 14306 17646 14306 17646 0 _371_
rlabel metal1 6992 16150 6992 16150 0 _372_
rlabel metal1 6118 18394 6118 18394 0 _373_
rlabel metal1 5796 18938 5796 18938 0 _374_
rlabel metal1 10166 17850 10166 17850 0 _375_
rlabel metal1 9200 18258 9200 18258 0 _376_
rlabel metal2 13754 18326 13754 18326 0 _377_
rlabel metal1 13432 17850 13432 17850 0 _378_
rlabel metal1 13524 16082 13524 16082 0 _379_
rlabel metal2 14214 16694 14214 16694 0 _380_
rlabel metal2 9062 19142 9062 19142 0 _381_
rlabel metal1 12328 17646 12328 17646 0 _382_
rlabel metal2 12374 18836 12374 18836 0 _383_
rlabel metal2 10902 19142 10902 19142 0 _384_
rlabel metal2 7958 17340 7958 17340 0 _385_
rlabel metal1 9246 17238 9246 17238 0 _386_
rlabel viali 11914 17169 11914 17169 0 _387_
rlabel metal1 11454 16694 11454 16694 0 _388_
rlabel metal1 11684 19822 11684 19822 0 _389_
rlabel metal1 9246 17714 9246 17714 0 _390_
rlabel metal1 8924 16558 8924 16558 0 _391_
rlabel metal1 9062 16422 9062 16422 0 _392_
rlabel metal2 12282 18564 12282 18564 0 _393_
rlabel metal2 11086 17510 11086 17510 0 _394_
rlabel metal2 12466 16252 12466 16252 0 _395_
rlabel via2 11638 16235 11638 16235 0 _396_
rlabel metal1 13202 16218 13202 16218 0 _397_
rlabel metal2 12052 19346 12052 19346 0 _398_
rlabel metal2 11270 12036 11270 12036 0 _399_
rlabel metal1 2714 12274 2714 12274 0 _400_
rlabel viali 18443 12206 18443 12206 0 _401_
rlabel metal1 18446 2958 18446 2958 0 _402_
rlabel metal1 12834 6766 12834 6766 0 _403_
rlabel metal1 12650 9996 12650 9996 0 _404_
rlabel metal2 19366 4114 19366 4114 0 _405_
rlabel metal1 13754 6290 13754 6290 0 _406_
rlabel metal1 21896 8466 21896 8466 0 _407_
rlabel metal1 20746 3434 20746 3434 0 _408_
rlabel metal1 18170 6766 18170 6766 0 _409_
rlabel metal1 22632 4590 22632 4590 0 _410_
rlabel metal3 751 1156 751 1156 0 clockp[0]
rlabel metal3 621 2516 621 2516 0 clockp[1]
rlabel metal2 1518 6018 1518 6018 0 clockp_buffer_in\[0\]
rlabel metal1 4600 20434 4600 20434 0 clockp_buffer_in\[1\]
rlabel metal1 13938 11118 13938 11118 0 dco
rlabel via1 5933 1938 5933 1938 0 div[0]
rlabel metal1 5060 1326 5060 1326 0 div[1]
rlabel metal1 3174 4658 3174 4658 0 div[2]
rlabel via1 3373 5678 3373 5678 0 div[3]
rlabel metal2 5014 8313 5014 8313 0 div[4]
rlabel metal3 1004 8772 1004 8772 0 div[5]
rlabel metal2 6210 9945 6210 9945 0 div[6]
rlabel metal2 1334 10829 1334 10829 0 div[7]
rlabel metal1 6302 1938 6302 1938 0 dll_control.accum\[0\]
rlabel metal1 5382 1836 5382 1836 0 dll_control.accum\[1\]
rlabel metal1 7038 4250 7038 4250 0 dll_control.accum\[2\]
rlabel metal1 3404 5134 3404 5134 0 dll_control.accum\[3\]
rlabel metal1 5336 7378 5336 7378 0 dll_control.accum\[4\]
rlabel metal1 5750 9010 5750 9010 0 dll_control.accum\[5\]
rlabel metal2 3266 9792 3266 9792 0 dll_control.accum\[6\]
rlabel metal1 5382 10574 5382 10574 0 dll_control.accum\[7\]
rlabel via1 4830 8466 4830 8466 0 dll_control.accum\[8\]
rlabel viali 7997 6324 7997 6324 0 dll_control.count0\[0\]
rlabel metal1 8878 2414 8878 2414 0 dll_control.count0\[1\]
rlabel metal1 7820 6358 7820 6358 0 dll_control.count0\[2\]
rlabel metal1 10166 5542 10166 5542 0 dll_control.count0\[3\]
rlabel metal2 6670 7140 6670 7140 0 dll_control.count0\[4\]
rlabel metal1 7176 8942 7176 8942 0 dll_control.count0\[5\]
rlabel metal1 14122 10540 14122 10540 0 dll_control.count1\[0\]
rlabel metal1 13616 10982 13616 10982 0 dll_control.count1\[1\]
rlabel metal2 9522 10302 9522 10302 0 dll_control.count1\[2\]
rlabel metal1 18262 11832 18262 11832 0 dll_control.count1\[3\]
rlabel metal2 18078 10880 18078 10880 0 dll_control.count1\[4\]
rlabel metal1 19136 9010 19136 9010 0 dll_control.count1\[5\]
rlabel metal1 15272 10098 15272 10098 0 dll_control.count2\[0\]
rlabel metal1 15916 10642 15916 10642 0 dll_control.count2\[1\]
rlabel metal2 16606 10914 16606 10914 0 dll_control.count2\[2\]
rlabel metal2 21022 11628 21022 11628 0 dll_control.count2\[3\]
rlabel metal1 21114 11594 21114 11594 0 dll_control.count2\[4\]
rlabel metal1 21390 9486 21390 9486 0 dll_control.count2\[5\]
rlabel metal2 15318 9418 15318 9418 0 dll_control.count3\[0\]
rlabel metal1 18584 10030 18584 10030 0 dll_control.count3\[1\]
rlabel metal1 18170 9486 18170 9486 0 dll_control.count3\[2\]
rlabel metal2 21942 8704 21942 8704 0 dll_control.count3\[3\]
rlabel metal1 23828 10438 23828 10438 0 dll_control.count3\[4\]
rlabel metal2 24794 9724 24794 9724 0 dll_control.count3\[5\]
rlabel metal1 14444 8398 14444 8398 0 dll_control.count4\[0\]
rlabel metal1 19734 4624 19734 4624 0 dll_control.count4\[1\]
rlabel metal1 17572 4250 17572 4250 0 dll_control.count4\[2\]
rlabel metal1 20930 6426 20930 6426 0 dll_control.count4\[3\]
rlabel metal1 24334 4454 24334 4454 0 dll_control.count4\[4\]
rlabel metal1 25024 6766 25024 6766 0 dll_control.count4\[5\]
rlabel metal2 14950 5984 14950 5984 0 dll_control.count5\[0\]
rlabel metal1 19872 4454 19872 4454 0 dll_control.count5\[1\]
rlabel metal1 17526 4046 17526 4046 0 dll_control.count5\[2\]
rlabel metal1 20746 5542 20746 5542 0 dll_control.count5\[3\]
rlabel metal1 23644 4998 23644 4998 0 dll_control.count5\[4\]
rlabel metal1 24334 6630 24334 6630 0 dll_control.count5\[5\]
rlabel metal1 15548 4454 15548 4454 0 dll_control.count6\[0\]
rlabel metal2 19734 1836 19734 1836 0 dll_control.count6\[1\]
rlabel metal1 16951 3094 16951 3094 0 dll_control.count6\[2\]
rlabel metal1 18216 5338 18216 5338 0 dll_control.count6\[3\]
rlabel metal1 22356 5338 22356 5338 0 dll_control.count6\[4\]
rlabel metal1 23874 6766 23874 6766 0 dll_control.count6\[5\]
rlabel metal2 13570 1530 13570 1530 0 dll_control.count7\[0\]
rlabel metal1 18078 2890 18078 2890 0 dll_control.count7\[1\]
rlabel metal1 13708 3366 13708 3366 0 dll_control.count7\[2\]
rlabel metal1 15180 5542 15180 5542 0 dll_control.count7\[3\]
rlabel metal1 22310 6222 22310 6222 0 dll_control.count7\[4\]
rlabel metal1 19320 9078 19320 9078 0 dll_control.count7\[5\]
rlabel metal1 12236 2074 12236 2074 0 dll_control.count8\[0\]
rlabel metal1 10764 3162 10764 3162 0 dll_control.count8\[1\]
rlabel metal1 8050 4556 8050 4556 0 dll_control.count8\[2\]
rlabel metal1 5290 4624 5290 4624 0 dll_control.count8\[3\]
rlabel metal2 11086 7072 11086 7072 0 dll_control.count8\[4\]
rlabel metal1 13110 8432 13110 8432 0 dll_control.count8\[5\]
rlabel metal2 21574 3264 21574 3264 0 dll_control.oscbuf\[0\]
rlabel metal1 19550 3570 19550 3570 0 dll_control.oscbuf\[1\]
rlabel metal1 16284 4726 16284 4726 0 dll_control.oscbuf\[2\]
rlabel metal1 9936 12886 9936 12886 0 dll_control.tint\[0\]
rlabel metal1 8832 15470 8832 15470 0 dll_control.tint\[1\]
rlabel metal2 12098 13668 12098 13668 0 dll_control.tint\[2\]
rlabel metal2 15870 14110 15870 14110 0 dll_control.tint\[3\]
rlabel metal1 15870 13498 15870 13498 0 dll_control.tint\[4\]
rlabel metal1 4186 14450 4186 14450 0 dll_control.tval\[0\]
rlabel metal2 3450 14314 3450 14314 0 dll_control.tval\[1\]
rlabel metal1 5106 14314 5106 14314 0 dll_control.tval\[2\]
rlabel metal3 1717 12036 1717 12036 0 enable
rlabel metal1 6624 18598 6624 18598 0 ext_trim[0]
rlabel metal2 15318 19584 15318 19584 0 ext_trim[10]
rlabel via1 14676 17646 14676 17646 0 ext_trim[11]
rlabel metal2 14122 19040 14122 19040 0 ext_trim[12]
rlabel metal2 13478 20648 13478 20648 0 ext_trim[13]
rlabel metal1 14306 19958 14306 19958 0 ext_trim[14]
rlabel metal2 13018 16048 13018 16048 0 ext_trim[15]
rlabel metal1 13018 17204 13018 17204 0 ext_trim[16]
rlabel metal2 21574 19118 21574 19118 0 ext_trim[17]
rlabel metal2 23598 19016 23598 19016 0 ext_trim[18]
rlabel metal2 25622 20274 25622 20274 0 ext_trim[19]
rlabel metal2 6946 17017 6946 17017 0 ext_trim[1]
rlabel metal2 24886 19805 24886 19805 0 ext_trim[20]
rlabel metal3 25630 16116 25630 16116 0 ext_trim[21]
rlabel metal3 25676 12580 25676 12580 0 ext_trim[22]
rlabel metal3 21168 9044 21168 9044 0 ext_trim[23]
rlabel metal3 26274 5508 26274 5508 0 ext_trim[24]
rlabel metal2 26312 1972 26312 1972 0 ext_trim[25]
rlabel metal2 7406 16473 7406 16473 0 ext_trim[2]
rlabel metal2 5658 17561 5658 17561 0 ext_trim[3]
rlabel metal2 4002 17561 4002 17561 0 ext_trim[4]
rlabel metal2 4646 19023 4646 19023 0 ext_trim[5]
rlabel metal1 6854 18190 6854 18190 0 ext_trim[6]
rlabel via1 1426 21301 1426 21301 0 ext_trim[7]
rlabel metal2 14582 19992 14582 19992 0 ext_trim[8]
rlabel metal2 5382 21226 5382 21226 0 ext_trim[9]
rlabel metal1 10718 12104 10718 12104 0 ireset
rlabel metal1 7452 19822 7452 19822 0 itrim\[0\]
rlabel metal1 16238 18258 16238 18258 0 itrim\[10\]
rlabel metal1 17342 17204 17342 17204 0 itrim\[11\]
rlabel metal1 14720 16150 14720 16150 0 itrim\[12\]
rlabel metal1 9246 19278 9246 19278 0 itrim\[13\]
rlabel metal2 10074 20128 10074 20128 0 itrim\[14\]
rlabel metal1 8418 17646 8418 17646 0 itrim\[15\]
rlabel metal1 8372 16014 8372 16014 0 itrim\[16\]
rlabel metal1 5106 17204 5106 17204 0 itrim\[17\]
rlabel metal2 5106 17986 5106 17986 0 itrim\[18\]
rlabel metal1 5014 19244 5014 19244 0 itrim\[19\]
rlabel metal1 8464 19346 8464 19346 0 itrim\[1\]
rlabel metal1 11500 20366 11500 20366 0 itrim\[20\]
rlabel metal1 14122 20366 14122 20366 0 itrim\[21\]
rlabel metal1 16146 19754 16146 19754 0 itrim\[22\]
rlabel metal1 16008 17850 16008 17850 0 itrim\[23\]
rlabel metal1 17158 16626 17158 16626 0 itrim\[24\]
rlabel metal2 16790 16524 16790 16524 0 itrim\[25\]
rlabel metal1 7452 16626 7452 16626 0 itrim\[2\]
rlabel metal1 5612 17170 5612 17170 0 itrim\[3\]
rlabel metal2 3910 16932 3910 16932 0 itrim\[4\]
rlabel metal1 4186 18190 4186 18190 0 itrim\[5\]
rlabel metal1 5290 19822 5290 19822 0 itrim\[6\]
rlabel metal2 13018 19108 13018 19108 0 itrim\[7\]
rlabel metal2 14214 19142 14214 19142 0 itrim\[8\]
rlabel metal1 15732 19278 15732 19278 0 itrim\[9\]
rlabel metal1 13800 16014 13800 16014 0 net104
rlabel metal1 13478 15572 13478 15572 0 net105
rlabel metal1 13156 14858 13156 14858 0 net106
rlabel metal2 13754 14790 13754 14790 0 net107
rlabel metal1 13018 14416 13018 14416 0 net108
rlabel metal1 15732 14586 15732 14586 0 net109
rlabel metal2 12650 14076 12650 14076 0 net110
rlabel metal1 9522 18836 9522 18836 0 net111
rlabel metal1 12742 14960 12742 14960 0 net112
rlabel metal2 4738 13056 4738 13056 0 net113
rlabel metal1 2714 15538 2714 15538 0 net114
rlabel metal1 2576 5678 2576 5678 0 net115
rlabel metal1 2162 7888 2162 7888 0 net116
rlabel metal2 9982 5440 9982 5440 0 net117
rlabel metal1 2576 15470 2576 15470 0 net118
rlabel metal1 8004 18802 8004 18802 0 net119
rlabel metal2 12466 18785 12466 18785 0 net120
rlabel metal1 14214 18360 14214 18360 0 net121
rlabel metal1 9062 16082 9062 16082 0 net122
rlabel metal2 9706 13141 9706 13141 0 net123
rlabel metal1 8694 14382 8694 14382 0 net124
rlabel metal2 9752 12580 9752 12580 0 net125
rlabel metal1 13018 4556 13018 4556 0 net126
rlabel metal1 12466 10064 12466 10064 0 net127
rlabel metal1 12218 7854 12218 7854 0 net128
rlabel metal1 14030 5202 14030 5202 0 net129
rlabel metal2 16698 3264 16698 3264 0 net130
rlabel metal2 23782 4590 23782 4590 0 net131
rlabel metal1 17940 6766 17940 6766 0 net132
rlabel via1 20102 7378 20102 7378 0 net133
rlabel metal1 18906 6290 18906 6290 0 net134
rlabel metal2 9154 16830 9154 16830 0 net135
rlabel metal1 9430 17680 9430 17680 0 net136
rlabel metal2 16192 16558 16192 16558 0 net137
rlabel metal1 17388 12410 17388 12410 0 net138
rlabel metal1 18354 6732 18354 6732 0 net139
rlabel metal2 20194 1095 20194 1095 0 osc
rlabel metal2 6762 959 6762 959 0 resetb
rlabel metal1 16928 14586 16928 14586 0 ringosc.c\[0\]
rlabel metal2 4830 19142 4830 19142 0 ringosc.c\[1\]
rlabel metal2 9430 20094 9430 20094 0 ringosc.dstage\[0\].id.d0
rlabel metal2 9430 19584 9430 19584 0 ringosc.dstage\[0\].id.d1
rlabel metal1 9062 19890 9062 19890 0 ringosc.dstage\[0\].id.d2
rlabel metal1 15870 16150 15870 16150 0 ringosc.dstage\[0\].id.in
rlabel metal1 8142 19958 8142 19958 0 ringosc.dstage\[0\].id.out
rlabel metal1 15502 17850 15502 17850 0 ringosc.dstage\[0\].id.ts
rlabel metal1 17158 17782 17158 17782 0 ringosc.dstage\[10\].id.d0
rlabel metal1 17296 17510 17296 17510 0 ringosc.dstage\[10\].id.d1
rlabel metal2 18170 18462 18170 18462 0 ringosc.dstage\[10\].id.d2
rlabel metal1 16422 19210 16422 19210 0 ringosc.dstage\[10\].id.in
rlabel metal1 17710 18122 17710 18122 0 ringosc.dstage\[10\].id.out
rlabel metal1 17342 18292 17342 18292 0 ringosc.dstage\[10\].id.ts
rlabel metal2 18446 17102 18446 17102 0 ringosc.dstage\[11\].id.d0
rlabel metal1 18124 16422 18124 16422 0 ringosc.dstage\[11\].id.d1
rlabel metal1 19136 16558 19136 16558 0 ringosc.dstage\[11\].id.d2
rlabel metal1 19090 17102 19090 17102 0 ringosc.dstage\[11\].id.out
rlabel metal2 18262 16864 18262 16864 0 ringosc.dstage\[11\].id.ts
rlabel metal1 10350 19924 10350 19924 0 ringosc.dstage\[1\].id.d0
rlabel viali 10178 20434 10178 20434 0 ringosc.dstage\[1\].id.d1
rlabel metal1 8280 19414 8280 19414 0 ringosc.dstage\[1\].id.d2
rlabel metal2 7498 19788 7498 19788 0 ringosc.dstage\[1\].id.out
rlabel metal1 10120 19822 10120 19822 0 ringosc.dstage\[1\].id.ts
rlabel metal1 8050 17782 8050 17782 0 ringosc.dstage\[2\].id.d0
rlabel metal1 7728 17510 7728 17510 0 ringosc.dstage\[2\].id.d1
rlabel metal1 6785 17102 6785 17102 0 ringosc.dstage\[2\].id.d2
rlabel metal2 7038 17442 7038 17442 0 ringosc.dstage\[2\].id.out
rlabel metal1 7590 17714 7590 17714 0 ringosc.dstage\[2\].id.ts
rlabel metal1 6992 15946 6992 15946 0 ringosc.dstage\[3\].id.d0
rlabel metal1 6486 16218 6486 16218 0 ringosc.dstage\[3\].id.d1
rlabel metal1 6371 15674 6371 15674 0 ringosc.dstage\[3\].id.d2
rlabel metal1 6072 16694 6072 16694 0 ringosc.dstage\[3\].id.out
rlabel metal1 6716 16082 6716 16082 0 ringosc.dstage\[3\].id.ts
rlabel metal1 4784 16762 4784 16762 0 ringosc.dstage\[4\].id.d0
rlabel metal1 4704 17646 4704 17646 0 ringosc.dstage\[4\].id.d1
rlabel metal2 4462 17374 4462 17374 0 ringosc.dstage\[4\].id.d2
rlabel metal2 4370 17408 4370 17408 0 ringosc.dstage\[4\].id.out
rlabel metal1 5152 16558 5152 16558 0 ringosc.dstage\[4\].id.ts
rlabel metal1 5612 18122 5612 18122 0 ringosc.dstage\[5\].id.d0
rlabel metal1 4002 18122 4002 18122 0 ringosc.dstage\[5\].id.d1
rlabel metal1 3703 18666 3703 18666 0 ringosc.dstage\[5\].id.d2
rlabel metal1 4048 18666 4048 18666 0 ringosc.dstage\[5\].id.out
rlabel metal1 4002 18258 4002 18258 0 ringosc.dstage\[5\].id.ts
rlabel metal1 5474 19278 5474 19278 0 ringosc.dstage\[6\].id.d0
rlabel metal1 5842 20570 5842 20570 0 ringosc.dstage\[6\].id.d1
rlabel metal1 5796 19890 5796 19890 0 ringosc.dstage\[6\].id.d2
rlabel metal1 5198 19958 5198 19958 0 ringosc.dstage\[6\].id.out
rlabel metal1 4876 19822 4876 19822 0 ringosc.dstage\[6\].id.ts
rlabel metal1 12144 20026 12144 20026 0 ringosc.dstage\[7\].id.d0
rlabel metal2 12742 19788 12742 19788 0 ringosc.dstage\[7\].id.d1
rlabel metal1 13501 19482 13501 19482 0 ringosc.dstage\[7\].id.d2
rlabel metal2 13754 20196 13754 20196 0 ringosc.dstage\[7\].id.out
rlabel metal2 12006 19924 12006 19924 0 ringosc.dstage\[7\].id.ts
rlabel metal2 14214 20162 14214 20162 0 ringosc.dstage\[8\].id.d0
rlabel metal1 15407 20434 15407 20434 0 ringosc.dstage\[8\].id.d1
rlabel metal2 15226 20060 15226 20060 0 ringosc.dstage\[8\].id.d2
rlabel metal1 15318 19754 15318 19754 0 ringosc.dstage\[8\].id.out
rlabel metal1 15502 19924 15502 19924 0 ringosc.dstage\[8\].id.ts
rlabel metal2 17250 20162 17250 20162 0 ringosc.dstage\[9\].id.d0
rlabel metal2 16330 20298 16330 20298 0 ringosc.dstage\[9\].id.d1
rlabel metal2 16790 19550 16790 19550 0 ringosc.dstage\[9\].id.d2
rlabel metal1 16974 19754 16974 19754 0 ringosc.dstage\[9\].id.ts
rlabel metal1 15364 16082 15364 16082 0 ringosc.iss.ctrl0
rlabel metal1 17296 15946 17296 15946 0 ringosc.iss.d0
rlabel metal2 16974 16932 16974 16932 0 ringosc.iss.d1
rlabel metal1 16560 15470 16560 15470 0 ringosc.iss.d2
rlabel metal2 16330 14722 16330 14722 0 ringosc.iss.one
<< properties >>
string FIXED_BBOX 0 0 27000 22000
<< end >>
