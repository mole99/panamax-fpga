VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO res_div
  CLASS BLOCK ;
  FOREIGN res_div ;
  ORIGIN 0.005 0.005 ;
  SIZE 20.680 BY 65.440 ;
  PIN vdda
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 0.605 62.740 1.915 64.845 ;
    END
  END vdda
  PIN vssa
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 18.755 62.740 20.065 64.845 ;
    END
  END vssa
  PIN vref
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 9.680 62.740 10.990 64.845 ;
    END
  END vref
  OBS
      LAYER pwell ;
        RECT -0.005 64.945 20.675 65.435 ;
        RECT -0.005 0.485 0.485 64.945 ;
        RECT 20.185 0.485 20.675 64.945 ;
        RECT -0.005 -0.005 20.675 0.485 ;
      LAYER li1 ;
        RECT 0.125 65.075 20.545 65.305 ;
        RECT 0.125 0.355 0.355 65.075 ;
        RECT 0.555 62.695 1.965 64.875 ;
        RECT 2.205 62.695 3.615 64.875 ;
        RECT 3.855 62.695 5.265 64.875 ;
        RECT 5.505 62.695 6.915 64.875 ;
        RECT 7.155 62.695 8.565 64.875 ;
        RECT 8.805 62.695 10.215 64.875 ;
        RECT 10.455 62.695 11.865 64.875 ;
        RECT 12.105 62.695 13.515 64.875 ;
        RECT 13.755 62.695 15.165 64.875 ;
        RECT 15.405 62.695 16.815 64.875 ;
        RECT 17.055 62.695 18.465 64.875 ;
        RECT 18.705 62.695 20.115 64.875 ;
        RECT 0.555 0.555 1.965 2.735 ;
        RECT 2.205 0.555 3.615 2.735 ;
        RECT 3.855 0.555 5.265 2.735 ;
        RECT 5.505 0.555 6.915 2.735 ;
        RECT 7.155 0.555 8.565 2.735 ;
        RECT 8.805 0.555 10.215 2.735 ;
        RECT 10.455 0.555 11.865 2.735 ;
        RECT 12.105 0.555 13.515 2.735 ;
        RECT 13.755 0.555 15.165 2.735 ;
        RECT 15.405 0.555 16.815 2.735 ;
        RECT 17.055 0.555 18.465 2.735 ;
        RECT 18.705 0.555 20.115 2.735 ;
        RECT 20.315 0.355 20.545 65.075 ;
        RECT 0.125 0.125 20.545 0.355 ;
      LAYER met1 ;
        RECT 0.125 65.075 20.545 65.305 ;
        RECT 0.125 0.355 0.355 65.075 ;
        RECT 0.605 62.740 1.915 64.845 ;
        RECT 2.255 62.740 5.215 64.845 ;
        RECT 5.555 62.740 8.515 64.845 ;
        RECT 8.855 62.740 11.815 64.845 ;
        RECT 12.155 62.740 15.115 64.845 ;
        RECT 15.455 62.740 18.415 64.845 ;
        RECT 18.755 62.740 20.545 65.075 ;
        RECT 0.605 0.585 3.565 2.690 ;
        RECT 3.905 0.585 6.865 2.690 ;
        RECT 7.205 0.585 10.165 2.690 ;
        RECT 10.505 0.585 13.465 2.690 ;
        RECT 13.805 0.585 16.765 2.690 ;
        RECT 17.105 0.585 20.065 2.690 ;
        RECT 20.315 0.355 20.545 62.740 ;
        RECT 0.125 0.125 20.545 0.355 ;
  END
END res_div
END LIBRARY

