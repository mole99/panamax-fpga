VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO follower_amp
  CLASS BLOCK ;
  FOREIGN follower_amp ;
  ORIGIN 0.130 7.610 ;
  SIZE 22.140 BY 63.375 ;
  PIN vsub
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -7.480 0.540 -6.735 ;
    END
  END vsub
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 1.380 52.410 2.380 53.410 ;
    END
  END vdd
  PIN out
    DIRECTION INOUT ;
    ANTENNAGATEAREA 2.400000 ;
    ANTENNADIFFAREA 48.430000 ;
    PORT
      LAYER met2 ;
        RECT 19.530 21.790 20.530 22.790 ;
    END
  END out
  PIN ena
    ANTENNAGATEAREA 0.702500 ;
    ANTENNADIFFAREA 0.202500 ;
    PORT
      LAYER met2 ;
        RECT 1.305 6.235 2.305 7.235 ;
    END
  END ena
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 1.415 9.875 2.415 10.875 ;
    END
  END vss
  PIN in
    DIRECTION INOUT ;
    ANTENNAGATEAREA 2.602500 ;
    ANTENNADIFFAREA 0.202500 ;
    PORT
      LAYER met2 ;
        RECT 1.285 14.900 2.285 15.900 ;
    END
  END in
  OBS
      LAYER pwell ;
        RECT -0.130 55.335 22.010 55.765 ;
        RECT -0.130 -7.180 0.300 55.335 ;
      LAYER nwell ;
        RECT 0.600 14.675 21.270 54.980 ;
        RECT 0.600 -5.300 2.175 14.675 ;
      LAYER pwell ;
        RECT 2.970 10.665 19.570 14.145 ;
        RECT 5.715 10.175 8.395 10.190 ;
        RECT 2.990 6.895 4.720 9.925 ;
        RECT 5.715 6.710 10.805 10.175 ;
        RECT 8.105 6.695 10.805 6.710 ;
        RECT 12.370 10.160 15.050 10.165 ;
        RECT 12.370 6.685 19.570 10.160 ;
        RECT 14.520 6.680 19.570 6.685 ;
        RECT 2.245 5.380 19.625 5.810 ;
        RECT 2.245 -4.800 2.675 5.380 ;
        RECT 19.195 -4.800 19.625 5.380 ;
        RECT 2.245 -5.230 19.625 -4.800 ;
      LAYER nwell ;
        RECT 19.695 -5.300 21.270 14.675 ;
        RECT 0.600 -6.875 21.270 -5.300 ;
      LAYER pwell ;
        RECT 21.580 -7.180 22.010 55.335 ;
        RECT -0.130 -7.610 22.010 -7.180 ;
      LAYER li1 ;
        RECT 0.000 55.145 21.885 55.645 ;
        RECT 0.000 -6.970 0.540 55.145 ;
        RECT 0.895 54.695 1.415 54.715 ;
        RECT 0.895 54.240 20.940 54.695 ;
        RECT 0.895 -6.075 1.415 54.240 ;
        RECT 1.860 53.215 19.865 53.660 ;
        RECT 1.860 22.360 2.710 53.215 ;
        RECT 3.295 52.660 3.795 52.830 ;
        RECT 4.085 52.660 4.585 52.830 ;
        RECT 4.875 52.660 5.375 52.830 ;
        RECT 5.665 52.660 6.165 52.830 ;
        RECT 6.455 52.660 6.955 52.830 ;
        RECT 7.245 52.660 7.745 52.830 ;
        RECT 8.035 52.660 8.535 52.830 ;
        RECT 8.825 52.660 9.325 52.830 ;
        RECT 9.615 52.660 10.115 52.830 ;
        RECT 10.405 52.660 10.905 52.830 ;
        RECT 11.195 52.660 11.695 52.830 ;
        RECT 11.985 52.660 12.485 52.830 ;
        RECT 12.775 52.660 13.275 52.830 ;
        RECT 13.565 52.660 14.065 52.830 ;
        RECT 14.355 52.660 14.855 52.830 ;
        RECT 15.145 52.660 15.645 52.830 ;
        RECT 15.935 52.660 16.435 52.830 ;
        RECT 16.725 52.660 17.225 52.830 ;
        RECT 17.515 52.660 18.015 52.830 ;
        RECT 18.305 52.660 18.805 52.830 ;
        RECT 3.065 51.405 3.235 52.445 ;
        RECT 3.855 51.405 4.025 52.445 ;
        RECT 4.645 51.405 4.815 52.445 ;
        RECT 5.435 51.405 5.605 52.445 ;
        RECT 6.225 51.405 6.395 52.445 ;
        RECT 7.015 51.405 7.185 52.445 ;
        RECT 7.805 51.405 7.975 52.445 ;
        RECT 8.595 51.405 8.765 52.445 ;
        RECT 9.385 51.405 9.555 52.445 ;
        RECT 10.175 51.405 10.345 52.445 ;
        RECT 10.965 51.405 11.135 52.445 ;
        RECT 11.755 51.405 11.925 52.445 ;
        RECT 12.545 51.405 12.715 52.445 ;
        RECT 13.335 51.405 13.505 52.445 ;
        RECT 14.125 51.405 14.295 52.445 ;
        RECT 14.915 51.405 15.085 52.445 ;
        RECT 15.705 51.405 15.875 52.445 ;
        RECT 16.495 51.405 16.665 52.445 ;
        RECT 17.285 51.405 17.455 52.445 ;
        RECT 18.075 51.405 18.245 52.445 ;
        RECT 18.865 51.405 19.035 52.445 ;
        RECT 3.295 51.020 3.795 51.190 ;
        RECT 4.085 51.020 4.585 51.190 ;
        RECT 4.875 51.020 5.375 51.190 ;
        RECT 5.665 51.020 6.165 51.190 ;
        RECT 6.455 51.020 6.955 51.190 ;
        RECT 7.245 51.020 7.745 51.190 ;
        RECT 8.035 51.020 8.535 51.190 ;
        RECT 8.825 51.020 9.325 51.190 ;
        RECT 9.615 51.020 10.115 51.190 ;
        RECT 10.405 51.020 10.905 51.190 ;
        RECT 11.195 51.020 11.695 51.190 ;
        RECT 11.985 51.020 12.485 51.190 ;
        RECT 12.775 51.020 13.275 51.190 ;
        RECT 13.565 51.020 14.065 51.190 ;
        RECT 14.355 51.020 14.855 51.190 ;
        RECT 15.145 51.020 15.645 51.190 ;
        RECT 15.935 51.020 16.435 51.190 ;
        RECT 16.725 51.020 17.225 51.190 ;
        RECT 17.515 51.020 18.015 51.190 ;
        RECT 18.305 51.020 18.805 51.190 ;
        RECT 3.295 50.480 3.795 50.650 ;
        RECT 4.085 50.480 4.585 50.650 ;
        RECT 4.875 50.480 5.375 50.650 ;
        RECT 5.665 50.480 6.165 50.650 ;
        RECT 6.455 50.480 6.955 50.650 ;
        RECT 7.245 50.480 7.745 50.650 ;
        RECT 8.035 50.480 8.535 50.650 ;
        RECT 8.825 50.480 9.325 50.650 ;
        RECT 9.615 50.480 10.115 50.650 ;
        RECT 10.405 50.480 10.905 50.650 ;
        RECT 11.195 50.480 11.695 50.650 ;
        RECT 11.985 50.480 12.485 50.650 ;
        RECT 12.775 50.480 13.275 50.650 ;
        RECT 13.565 50.480 14.065 50.650 ;
        RECT 14.355 50.480 14.855 50.650 ;
        RECT 15.145 50.480 15.645 50.650 ;
        RECT 15.935 50.480 16.435 50.650 ;
        RECT 16.725 50.480 17.225 50.650 ;
        RECT 17.515 50.480 18.015 50.650 ;
        RECT 18.305 50.480 18.805 50.650 ;
        RECT 3.065 49.225 3.235 50.265 ;
        RECT 3.855 49.225 4.025 50.265 ;
        RECT 4.645 49.225 4.815 50.265 ;
        RECT 5.435 49.225 5.605 50.265 ;
        RECT 6.225 49.225 6.395 50.265 ;
        RECT 7.015 49.225 7.185 50.265 ;
        RECT 7.805 49.225 7.975 50.265 ;
        RECT 8.595 49.225 8.765 50.265 ;
        RECT 9.385 49.225 9.555 50.265 ;
        RECT 10.175 49.225 10.345 50.265 ;
        RECT 10.965 49.225 11.135 50.265 ;
        RECT 11.755 49.225 11.925 50.265 ;
        RECT 12.545 49.225 12.715 50.265 ;
        RECT 13.335 49.225 13.505 50.265 ;
        RECT 14.125 49.225 14.295 50.265 ;
        RECT 14.915 49.225 15.085 50.265 ;
        RECT 15.705 49.225 15.875 50.265 ;
        RECT 16.495 49.225 16.665 50.265 ;
        RECT 17.285 49.225 17.455 50.265 ;
        RECT 18.075 49.225 18.245 50.265 ;
        RECT 18.865 49.225 19.035 50.265 ;
        RECT 3.295 48.840 3.795 49.010 ;
        RECT 4.085 48.840 4.585 49.010 ;
        RECT 4.875 48.840 5.375 49.010 ;
        RECT 5.665 48.840 6.165 49.010 ;
        RECT 6.455 48.840 6.955 49.010 ;
        RECT 7.245 48.840 7.745 49.010 ;
        RECT 8.035 48.840 8.535 49.010 ;
        RECT 8.825 48.840 9.325 49.010 ;
        RECT 9.615 48.840 10.115 49.010 ;
        RECT 10.405 48.840 10.905 49.010 ;
        RECT 11.195 48.840 11.695 49.010 ;
        RECT 11.985 48.840 12.485 49.010 ;
        RECT 12.775 48.840 13.275 49.010 ;
        RECT 13.565 48.840 14.065 49.010 ;
        RECT 14.355 48.840 14.855 49.010 ;
        RECT 15.145 48.840 15.645 49.010 ;
        RECT 15.935 48.840 16.435 49.010 ;
        RECT 16.725 48.840 17.225 49.010 ;
        RECT 17.515 48.840 18.015 49.010 ;
        RECT 18.305 48.840 18.805 49.010 ;
        RECT 3.295 48.300 3.795 48.470 ;
        RECT 4.085 48.300 4.585 48.470 ;
        RECT 4.875 48.300 5.375 48.470 ;
        RECT 5.665 48.300 6.165 48.470 ;
        RECT 6.455 48.300 6.955 48.470 ;
        RECT 7.245 48.300 7.745 48.470 ;
        RECT 8.035 48.300 8.535 48.470 ;
        RECT 8.825 48.300 9.325 48.470 ;
        RECT 9.615 48.300 10.115 48.470 ;
        RECT 10.405 48.300 10.905 48.470 ;
        RECT 11.195 48.300 11.695 48.470 ;
        RECT 11.985 48.300 12.485 48.470 ;
        RECT 12.775 48.300 13.275 48.470 ;
        RECT 13.565 48.300 14.065 48.470 ;
        RECT 14.355 48.300 14.855 48.470 ;
        RECT 15.145 48.300 15.645 48.470 ;
        RECT 15.935 48.300 16.435 48.470 ;
        RECT 16.725 48.300 17.225 48.470 ;
        RECT 17.515 48.300 18.015 48.470 ;
        RECT 18.305 48.300 18.805 48.470 ;
        RECT 3.065 47.045 3.235 48.085 ;
        RECT 3.855 47.045 4.025 48.085 ;
        RECT 4.645 47.045 4.815 48.085 ;
        RECT 5.435 47.045 5.605 48.085 ;
        RECT 6.225 47.045 6.395 48.085 ;
        RECT 7.015 47.045 7.185 48.085 ;
        RECT 7.805 47.045 7.975 48.085 ;
        RECT 8.595 47.045 8.765 48.085 ;
        RECT 9.385 47.045 9.555 48.085 ;
        RECT 10.175 47.045 10.345 48.085 ;
        RECT 10.965 47.045 11.135 48.085 ;
        RECT 11.755 47.045 11.925 48.085 ;
        RECT 12.545 47.045 12.715 48.085 ;
        RECT 13.335 47.045 13.505 48.085 ;
        RECT 14.125 47.045 14.295 48.085 ;
        RECT 14.915 47.045 15.085 48.085 ;
        RECT 15.705 47.045 15.875 48.085 ;
        RECT 16.495 47.045 16.665 48.085 ;
        RECT 17.285 47.045 17.455 48.085 ;
        RECT 18.075 47.045 18.245 48.085 ;
        RECT 18.865 47.045 19.035 48.085 ;
        RECT 3.295 46.660 3.795 46.830 ;
        RECT 4.085 46.660 4.585 46.830 ;
        RECT 4.875 46.660 5.375 46.830 ;
        RECT 5.665 46.660 6.165 46.830 ;
        RECT 6.455 46.660 6.955 46.830 ;
        RECT 7.245 46.660 7.745 46.830 ;
        RECT 8.035 46.660 8.535 46.830 ;
        RECT 8.825 46.660 9.325 46.830 ;
        RECT 9.615 46.660 10.115 46.830 ;
        RECT 10.405 46.660 10.905 46.830 ;
        RECT 11.195 46.660 11.695 46.830 ;
        RECT 11.985 46.660 12.485 46.830 ;
        RECT 12.775 46.660 13.275 46.830 ;
        RECT 13.565 46.660 14.065 46.830 ;
        RECT 14.355 46.660 14.855 46.830 ;
        RECT 15.145 46.660 15.645 46.830 ;
        RECT 15.935 46.660 16.435 46.830 ;
        RECT 16.725 46.660 17.225 46.830 ;
        RECT 17.515 46.660 18.015 46.830 ;
        RECT 18.305 46.660 18.805 46.830 ;
        RECT 3.295 46.120 3.795 46.290 ;
        RECT 4.085 46.120 4.585 46.290 ;
        RECT 4.875 46.120 5.375 46.290 ;
        RECT 5.665 46.120 6.165 46.290 ;
        RECT 6.455 46.120 6.955 46.290 ;
        RECT 7.245 46.120 7.745 46.290 ;
        RECT 8.035 46.120 8.535 46.290 ;
        RECT 8.825 46.120 9.325 46.290 ;
        RECT 9.615 46.120 10.115 46.290 ;
        RECT 10.405 46.120 10.905 46.290 ;
        RECT 11.195 46.120 11.695 46.290 ;
        RECT 11.985 46.120 12.485 46.290 ;
        RECT 12.775 46.120 13.275 46.290 ;
        RECT 13.565 46.120 14.065 46.290 ;
        RECT 14.355 46.120 14.855 46.290 ;
        RECT 15.145 46.120 15.645 46.290 ;
        RECT 15.935 46.120 16.435 46.290 ;
        RECT 16.725 46.120 17.225 46.290 ;
        RECT 17.515 46.120 18.015 46.290 ;
        RECT 18.305 46.120 18.805 46.290 ;
        RECT 3.065 44.865 3.235 45.905 ;
        RECT 3.855 44.865 4.025 45.905 ;
        RECT 4.645 44.865 4.815 45.905 ;
        RECT 5.435 44.865 5.605 45.905 ;
        RECT 6.225 44.865 6.395 45.905 ;
        RECT 7.015 44.865 7.185 45.905 ;
        RECT 7.805 44.865 7.975 45.905 ;
        RECT 8.595 44.865 8.765 45.905 ;
        RECT 9.385 44.865 9.555 45.905 ;
        RECT 10.175 44.865 10.345 45.905 ;
        RECT 10.965 44.865 11.135 45.905 ;
        RECT 11.755 44.865 11.925 45.905 ;
        RECT 12.545 44.865 12.715 45.905 ;
        RECT 13.335 44.865 13.505 45.905 ;
        RECT 14.125 44.865 14.295 45.905 ;
        RECT 14.915 44.865 15.085 45.905 ;
        RECT 15.705 44.865 15.875 45.905 ;
        RECT 16.495 44.865 16.665 45.905 ;
        RECT 17.285 44.865 17.455 45.905 ;
        RECT 18.075 44.865 18.245 45.905 ;
        RECT 18.865 44.865 19.035 45.905 ;
        RECT 3.295 44.480 3.795 44.650 ;
        RECT 4.085 44.480 4.585 44.650 ;
        RECT 4.875 44.480 5.375 44.650 ;
        RECT 5.665 44.480 6.165 44.650 ;
        RECT 6.455 44.480 6.955 44.650 ;
        RECT 7.245 44.480 7.745 44.650 ;
        RECT 8.035 44.480 8.535 44.650 ;
        RECT 8.825 44.480 9.325 44.650 ;
        RECT 9.615 44.480 10.115 44.650 ;
        RECT 10.405 44.480 10.905 44.650 ;
        RECT 11.195 44.480 11.695 44.650 ;
        RECT 11.985 44.480 12.485 44.650 ;
        RECT 12.775 44.480 13.275 44.650 ;
        RECT 13.565 44.480 14.065 44.650 ;
        RECT 14.355 44.480 14.855 44.650 ;
        RECT 15.145 44.480 15.645 44.650 ;
        RECT 15.935 44.480 16.435 44.650 ;
        RECT 16.725 44.480 17.225 44.650 ;
        RECT 17.515 44.480 18.015 44.650 ;
        RECT 18.305 44.480 18.805 44.650 ;
        RECT 3.295 43.940 3.795 44.110 ;
        RECT 4.085 43.940 4.585 44.110 ;
        RECT 4.875 43.940 5.375 44.110 ;
        RECT 5.665 43.940 6.165 44.110 ;
        RECT 6.455 43.940 6.955 44.110 ;
        RECT 7.245 43.940 7.745 44.110 ;
        RECT 8.035 43.940 8.535 44.110 ;
        RECT 8.825 43.940 9.325 44.110 ;
        RECT 9.615 43.940 10.115 44.110 ;
        RECT 10.405 43.940 10.905 44.110 ;
        RECT 11.195 43.940 11.695 44.110 ;
        RECT 11.985 43.940 12.485 44.110 ;
        RECT 12.775 43.940 13.275 44.110 ;
        RECT 13.565 43.940 14.065 44.110 ;
        RECT 14.355 43.940 14.855 44.110 ;
        RECT 15.145 43.940 15.645 44.110 ;
        RECT 15.935 43.940 16.435 44.110 ;
        RECT 16.725 43.940 17.225 44.110 ;
        RECT 17.515 43.940 18.015 44.110 ;
        RECT 18.305 43.940 18.805 44.110 ;
        RECT 3.065 42.685 3.235 43.725 ;
        RECT 3.855 42.685 4.025 43.725 ;
        RECT 4.645 42.685 4.815 43.725 ;
        RECT 5.435 42.685 5.605 43.725 ;
        RECT 6.225 42.685 6.395 43.725 ;
        RECT 7.015 42.685 7.185 43.725 ;
        RECT 7.805 42.685 7.975 43.725 ;
        RECT 8.595 42.685 8.765 43.725 ;
        RECT 9.385 42.685 9.555 43.725 ;
        RECT 10.175 42.685 10.345 43.725 ;
        RECT 10.965 42.685 11.135 43.725 ;
        RECT 11.755 42.685 11.925 43.725 ;
        RECT 12.545 42.685 12.715 43.725 ;
        RECT 13.335 42.685 13.505 43.725 ;
        RECT 14.125 42.685 14.295 43.725 ;
        RECT 14.915 42.685 15.085 43.725 ;
        RECT 15.705 42.685 15.875 43.725 ;
        RECT 16.495 42.685 16.665 43.725 ;
        RECT 17.285 42.685 17.455 43.725 ;
        RECT 18.075 42.685 18.245 43.725 ;
        RECT 18.865 42.685 19.035 43.725 ;
        RECT 3.295 42.300 3.795 42.470 ;
        RECT 4.085 42.300 4.585 42.470 ;
        RECT 4.875 42.300 5.375 42.470 ;
        RECT 5.665 42.300 6.165 42.470 ;
        RECT 6.455 42.300 6.955 42.470 ;
        RECT 7.245 42.300 7.745 42.470 ;
        RECT 8.035 42.300 8.535 42.470 ;
        RECT 8.825 42.300 9.325 42.470 ;
        RECT 9.615 42.300 10.115 42.470 ;
        RECT 10.405 42.300 10.905 42.470 ;
        RECT 11.195 42.300 11.695 42.470 ;
        RECT 11.985 42.300 12.485 42.470 ;
        RECT 12.775 42.300 13.275 42.470 ;
        RECT 13.565 42.300 14.065 42.470 ;
        RECT 14.355 42.300 14.855 42.470 ;
        RECT 15.145 42.300 15.645 42.470 ;
        RECT 15.935 42.300 16.435 42.470 ;
        RECT 16.725 42.300 17.225 42.470 ;
        RECT 17.515 42.300 18.015 42.470 ;
        RECT 18.305 42.300 18.805 42.470 ;
        RECT 3.295 41.760 3.795 41.930 ;
        RECT 4.085 41.760 4.585 41.930 ;
        RECT 4.875 41.760 5.375 41.930 ;
        RECT 5.665 41.760 6.165 41.930 ;
        RECT 6.455 41.760 6.955 41.930 ;
        RECT 7.245 41.760 7.745 41.930 ;
        RECT 8.035 41.760 8.535 41.930 ;
        RECT 8.825 41.760 9.325 41.930 ;
        RECT 9.615 41.760 10.115 41.930 ;
        RECT 10.405 41.760 10.905 41.930 ;
        RECT 11.195 41.760 11.695 41.930 ;
        RECT 11.985 41.760 12.485 41.930 ;
        RECT 12.775 41.760 13.275 41.930 ;
        RECT 13.565 41.760 14.065 41.930 ;
        RECT 14.355 41.760 14.855 41.930 ;
        RECT 15.145 41.760 15.645 41.930 ;
        RECT 15.935 41.760 16.435 41.930 ;
        RECT 16.725 41.760 17.225 41.930 ;
        RECT 17.515 41.760 18.015 41.930 ;
        RECT 18.305 41.760 18.805 41.930 ;
        RECT 3.065 40.505 3.235 41.545 ;
        RECT 3.855 40.505 4.025 41.545 ;
        RECT 4.645 40.505 4.815 41.545 ;
        RECT 5.435 40.505 5.605 41.545 ;
        RECT 6.225 40.505 6.395 41.545 ;
        RECT 7.015 40.505 7.185 41.545 ;
        RECT 7.805 40.505 7.975 41.545 ;
        RECT 8.595 40.505 8.765 41.545 ;
        RECT 9.385 40.505 9.555 41.545 ;
        RECT 10.175 40.505 10.345 41.545 ;
        RECT 10.965 40.505 11.135 41.545 ;
        RECT 11.755 40.505 11.925 41.545 ;
        RECT 12.545 40.505 12.715 41.545 ;
        RECT 13.335 40.505 13.505 41.545 ;
        RECT 14.125 40.505 14.295 41.545 ;
        RECT 14.915 40.505 15.085 41.545 ;
        RECT 15.705 40.505 15.875 41.545 ;
        RECT 16.495 40.505 16.665 41.545 ;
        RECT 17.285 40.505 17.455 41.545 ;
        RECT 18.075 40.505 18.245 41.545 ;
        RECT 18.865 40.505 19.035 41.545 ;
        RECT 3.295 40.120 3.795 40.290 ;
        RECT 4.085 40.120 4.585 40.290 ;
        RECT 4.875 40.120 5.375 40.290 ;
        RECT 5.665 40.120 6.165 40.290 ;
        RECT 6.455 40.120 6.955 40.290 ;
        RECT 7.245 40.120 7.745 40.290 ;
        RECT 8.035 40.120 8.535 40.290 ;
        RECT 8.825 40.120 9.325 40.290 ;
        RECT 9.615 40.120 10.115 40.290 ;
        RECT 10.405 40.120 10.905 40.290 ;
        RECT 11.195 40.120 11.695 40.290 ;
        RECT 11.985 40.120 12.485 40.290 ;
        RECT 12.775 40.120 13.275 40.290 ;
        RECT 13.565 40.120 14.065 40.290 ;
        RECT 14.355 40.120 14.855 40.290 ;
        RECT 15.145 40.120 15.645 40.290 ;
        RECT 15.935 40.120 16.435 40.290 ;
        RECT 16.725 40.120 17.225 40.290 ;
        RECT 17.515 40.120 18.015 40.290 ;
        RECT 18.305 40.120 18.805 40.290 ;
        RECT 3.295 39.580 3.795 39.750 ;
        RECT 4.085 39.580 4.585 39.750 ;
        RECT 4.875 39.580 5.375 39.750 ;
        RECT 5.665 39.580 6.165 39.750 ;
        RECT 6.455 39.580 6.955 39.750 ;
        RECT 7.245 39.580 7.745 39.750 ;
        RECT 8.035 39.580 8.535 39.750 ;
        RECT 8.825 39.580 9.325 39.750 ;
        RECT 9.615 39.580 10.115 39.750 ;
        RECT 10.405 39.580 10.905 39.750 ;
        RECT 11.195 39.580 11.695 39.750 ;
        RECT 11.985 39.580 12.485 39.750 ;
        RECT 12.775 39.580 13.275 39.750 ;
        RECT 13.565 39.580 14.065 39.750 ;
        RECT 14.355 39.580 14.855 39.750 ;
        RECT 15.145 39.580 15.645 39.750 ;
        RECT 15.935 39.580 16.435 39.750 ;
        RECT 16.725 39.580 17.225 39.750 ;
        RECT 17.515 39.580 18.015 39.750 ;
        RECT 18.305 39.580 18.805 39.750 ;
        RECT 3.065 38.325 3.235 39.365 ;
        RECT 3.855 38.325 4.025 39.365 ;
        RECT 4.645 38.325 4.815 39.365 ;
        RECT 5.435 38.325 5.605 39.365 ;
        RECT 6.225 38.325 6.395 39.365 ;
        RECT 7.015 38.325 7.185 39.365 ;
        RECT 7.805 38.325 7.975 39.365 ;
        RECT 8.595 38.325 8.765 39.365 ;
        RECT 9.385 38.325 9.555 39.365 ;
        RECT 10.175 38.325 10.345 39.365 ;
        RECT 10.965 38.325 11.135 39.365 ;
        RECT 11.755 38.325 11.925 39.365 ;
        RECT 12.545 38.325 12.715 39.365 ;
        RECT 13.335 38.325 13.505 39.365 ;
        RECT 14.125 38.325 14.295 39.365 ;
        RECT 14.915 38.325 15.085 39.365 ;
        RECT 15.705 38.325 15.875 39.365 ;
        RECT 16.495 38.325 16.665 39.365 ;
        RECT 17.285 38.325 17.455 39.365 ;
        RECT 18.075 38.325 18.245 39.365 ;
        RECT 18.865 38.325 19.035 39.365 ;
        RECT 3.295 37.940 3.795 38.110 ;
        RECT 4.085 37.940 4.585 38.110 ;
        RECT 4.875 37.940 5.375 38.110 ;
        RECT 5.665 37.940 6.165 38.110 ;
        RECT 6.455 37.940 6.955 38.110 ;
        RECT 7.245 37.940 7.745 38.110 ;
        RECT 8.035 37.940 8.535 38.110 ;
        RECT 8.825 37.940 9.325 38.110 ;
        RECT 9.615 37.940 10.115 38.110 ;
        RECT 10.405 37.940 10.905 38.110 ;
        RECT 11.195 37.940 11.695 38.110 ;
        RECT 11.985 37.940 12.485 38.110 ;
        RECT 12.775 37.940 13.275 38.110 ;
        RECT 13.565 37.940 14.065 38.110 ;
        RECT 14.355 37.940 14.855 38.110 ;
        RECT 15.145 37.940 15.645 38.110 ;
        RECT 15.935 37.940 16.435 38.110 ;
        RECT 16.725 37.940 17.225 38.110 ;
        RECT 17.515 37.940 18.015 38.110 ;
        RECT 18.305 37.940 18.805 38.110 ;
        RECT 3.295 37.400 3.795 37.570 ;
        RECT 4.085 37.400 4.585 37.570 ;
        RECT 4.875 37.400 5.375 37.570 ;
        RECT 5.665 37.400 6.165 37.570 ;
        RECT 6.455 37.400 6.955 37.570 ;
        RECT 7.245 37.400 7.745 37.570 ;
        RECT 8.035 37.400 8.535 37.570 ;
        RECT 8.825 37.400 9.325 37.570 ;
        RECT 9.615 37.400 10.115 37.570 ;
        RECT 10.405 37.400 10.905 37.570 ;
        RECT 11.195 37.400 11.695 37.570 ;
        RECT 11.985 37.400 12.485 37.570 ;
        RECT 12.775 37.400 13.275 37.570 ;
        RECT 13.565 37.400 14.065 37.570 ;
        RECT 14.355 37.400 14.855 37.570 ;
        RECT 15.145 37.400 15.645 37.570 ;
        RECT 15.935 37.400 16.435 37.570 ;
        RECT 16.725 37.400 17.225 37.570 ;
        RECT 17.515 37.400 18.015 37.570 ;
        RECT 18.305 37.400 18.805 37.570 ;
        RECT 3.065 36.145 3.235 37.185 ;
        RECT 3.855 36.145 4.025 37.185 ;
        RECT 4.645 36.145 4.815 37.185 ;
        RECT 5.435 36.145 5.605 37.185 ;
        RECT 6.225 36.145 6.395 37.185 ;
        RECT 7.015 36.145 7.185 37.185 ;
        RECT 7.805 36.145 7.975 37.185 ;
        RECT 8.595 36.145 8.765 37.185 ;
        RECT 9.385 36.145 9.555 37.185 ;
        RECT 10.175 36.145 10.345 37.185 ;
        RECT 10.965 36.145 11.135 37.185 ;
        RECT 11.755 36.145 11.925 37.185 ;
        RECT 12.545 36.145 12.715 37.185 ;
        RECT 13.335 36.145 13.505 37.185 ;
        RECT 14.125 36.145 14.295 37.185 ;
        RECT 14.915 36.145 15.085 37.185 ;
        RECT 15.705 36.145 15.875 37.185 ;
        RECT 16.495 36.145 16.665 37.185 ;
        RECT 17.285 36.145 17.455 37.185 ;
        RECT 18.075 36.145 18.245 37.185 ;
        RECT 18.865 36.145 19.035 37.185 ;
        RECT 3.295 35.760 3.795 35.930 ;
        RECT 4.085 35.760 4.585 35.930 ;
        RECT 4.875 35.760 5.375 35.930 ;
        RECT 5.665 35.760 6.165 35.930 ;
        RECT 6.455 35.760 6.955 35.930 ;
        RECT 7.245 35.760 7.745 35.930 ;
        RECT 8.035 35.760 8.535 35.930 ;
        RECT 8.825 35.760 9.325 35.930 ;
        RECT 9.615 35.760 10.115 35.930 ;
        RECT 10.405 35.760 10.905 35.930 ;
        RECT 11.195 35.760 11.695 35.930 ;
        RECT 11.985 35.760 12.485 35.930 ;
        RECT 12.775 35.760 13.275 35.930 ;
        RECT 13.565 35.760 14.065 35.930 ;
        RECT 14.355 35.760 14.855 35.930 ;
        RECT 15.145 35.760 15.645 35.930 ;
        RECT 15.935 35.760 16.435 35.930 ;
        RECT 16.725 35.760 17.225 35.930 ;
        RECT 17.515 35.760 18.015 35.930 ;
        RECT 18.305 35.760 18.805 35.930 ;
        RECT 3.295 35.220 3.795 35.390 ;
        RECT 4.085 35.220 4.585 35.390 ;
        RECT 4.875 35.220 5.375 35.390 ;
        RECT 5.665 35.220 6.165 35.390 ;
        RECT 6.455 35.220 6.955 35.390 ;
        RECT 7.245 35.220 7.745 35.390 ;
        RECT 8.035 35.220 8.535 35.390 ;
        RECT 8.825 35.220 9.325 35.390 ;
        RECT 9.615 35.220 10.115 35.390 ;
        RECT 10.405 35.220 10.905 35.390 ;
        RECT 11.195 35.220 11.695 35.390 ;
        RECT 11.985 35.220 12.485 35.390 ;
        RECT 12.775 35.220 13.275 35.390 ;
        RECT 13.565 35.220 14.065 35.390 ;
        RECT 14.355 35.220 14.855 35.390 ;
        RECT 15.145 35.220 15.645 35.390 ;
        RECT 15.935 35.220 16.435 35.390 ;
        RECT 16.725 35.220 17.225 35.390 ;
        RECT 17.515 35.220 18.015 35.390 ;
        RECT 18.305 35.220 18.805 35.390 ;
        RECT 3.065 33.965 3.235 35.005 ;
        RECT 3.855 33.965 4.025 35.005 ;
        RECT 4.645 33.965 4.815 35.005 ;
        RECT 5.435 33.965 5.605 35.005 ;
        RECT 6.225 33.965 6.395 35.005 ;
        RECT 7.015 33.965 7.185 35.005 ;
        RECT 7.805 33.965 7.975 35.005 ;
        RECT 8.595 33.965 8.765 35.005 ;
        RECT 9.385 33.965 9.555 35.005 ;
        RECT 10.175 33.965 10.345 35.005 ;
        RECT 10.965 33.965 11.135 35.005 ;
        RECT 11.755 33.965 11.925 35.005 ;
        RECT 12.545 33.965 12.715 35.005 ;
        RECT 13.335 33.965 13.505 35.005 ;
        RECT 14.125 33.965 14.295 35.005 ;
        RECT 14.915 33.965 15.085 35.005 ;
        RECT 15.705 33.965 15.875 35.005 ;
        RECT 16.495 33.965 16.665 35.005 ;
        RECT 17.285 33.965 17.455 35.005 ;
        RECT 18.075 33.965 18.245 35.005 ;
        RECT 18.865 33.965 19.035 35.005 ;
        RECT 3.295 33.580 3.795 33.750 ;
        RECT 4.085 33.580 4.585 33.750 ;
        RECT 4.875 33.580 5.375 33.750 ;
        RECT 5.665 33.580 6.165 33.750 ;
        RECT 6.455 33.580 6.955 33.750 ;
        RECT 7.245 33.580 7.745 33.750 ;
        RECT 8.035 33.580 8.535 33.750 ;
        RECT 8.825 33.580 9.325 33.750 ;
        RECT 9.615 33.580 10.115 33.750 ;
        RECT 10.405 33.580 10.905 33.750 ;
        RECT 11.195 33.580 11.695 33.750 ;
        RECT 11.985 33.580 12.485 33.750 ;
        RECT 12.775 33.580 13.275 33.750 ;
        RECT 13.565 33.580 14.065 33.750 ;
        RECT 14.355 33.580 14.855 33.750 ;
        RECT 15.145 33.580 15.645 33.750 ;
        RECT 15.935 33.580 16.435 33.750 ;
        RECT 16.725 33.580 17.225 33.750 ;
        RECT 17.515 33.580 18.015 33.750 ;
        RECT 18.305 33.580 18.805 33.750 ;
        RECT 3.295 33.040 3.795 33.210 ;
        RECT 4.085 33.040 4.585 33.210 ;
        RECT 4.875 33.040 5.375 33.210 ;
        RECT 5.665 33.040 6.165 33.210 ;
        RECT 6.455 33.040 6.955 33.210 ;
        RECT 7.245 33.040 7.745 33.210 ;
        RECT 8.035 33.040 8.535 33.210 ;
        RECT 8.825 33.040 9.325 33.210 ;
        RECT 9.615 33.040 10.115 33.210 ;
        RECT 10.405 33.040 10.905 33.210 ;
        RECT 11.195 33.040 11.695 33.210 ;
        RECT 11.985 33.040 12.485 33.210 ;
        RECT 12.775 33.040 13.275 33.210 ;
        RECT 13.565 33.040 14.065 33.210 ;
        RECT 14.355 33.040 14.855 33.210 ;
        RECT 15.145 33.040 15.645 33.210 ;
        RECT 15.935 33.040 16.435 33.210 ;
        RECT 16.725 33.040 17.225 33.210 ;
        RECT 17.515 33.040 18.015 33.210 ;
        RECT 18.305 33.040 18.805 33.210 ;
        RECT 3.065 31.785 3.235 32.825 ;
        RECT 3.855 31.785 4.025 32.825 ;
        RECT 4.645 31.785 4.815 32.825 ;
        RECT 5.435 31.785 5.605 32.825 ;
        RECT 6.225 31.785 6.395 32.825 ;
        RECT 7.015 31.785 7.185 32.825 ;
        RECT 7.805 31.785 7.975 32.825 ;
        RECT 8.595 31.785 8.765 32.825 ;
        RECT 9.385 31.785 9.555 32.825 ;
        RECT 10.175 31.785 10.345 32.825 ;
        RECT 10.965 31.785 11.135 32.825 ;
        RECT 11.755 31.785 11.925 32.825 ;
        RECT 12.545 31.785 12.715 32.825 ;
        RECT 13.335 31.785 13.505 32.825 ;
        RECT 14.125 31.785 14.295 32.825 ;
        RECT 14.915 31.785 15.085 32.825 ;
        RECT 15.705 31.785 15.875 32.825 ;
        RECT 16.495 31.785 16.665 32.825 ;
        RECT 17.285 31.785 17.455 32.825 ;
        RECT 18.075 31.785 18.245 32.825 ;
        RECT 18.865 31.785 19.035 32.825 ;
        RECT 3.295 31.400 3.795 31.570 ;
        RECT 4.085 31.400 4.585 31.570 ;
        RECT 4.875 31.400 5.375 31.570 ;
        RECT 5.665 31.400 6.165 31.570 ;
        RECT 6.455 31.400 6.955 31.570 ;
        RECT 7.245 31.400 7.745 31.570 ;
        RECT 8.035 31.400 8.535 31.570 ;
        RECT 8.825 31.400 9.325 31.570 ;
        RECT 9.615 31.400 10.115 31.570 ;
        RECT 10.405 31.400 10.905 31.570 ;
        RECT 11.195 31.400 11.695 31.570 ;
        RECT 11.985 31.400 12.485 31.570 ;
        RECT 12.775 31.400 13.275 31.570 ;
        RECT 13.565 31.400 14.065 31.570 ;
        RECT 14.355 31.400 14.855 31.570 ;
        RECT 15.145 31.400 15.645 31.570 ;
        RECT 15.935 31.400 16.435 31.570 ;
        RECT 16.725 31.400 17.225 31.570 ;
        RECT 17.515 31.400 18.015 31.570 ;
        RECT 18.305 31.400 18.805 31.570 ;
        RECT 3.295 30.860 3.795 31.030 ;
        RECT 4.085 30.860 4.585 31.030 ;
        RECT 4.875 30.860 5.375 31.030 ;
        RECT 5.665 30.860 6.165 31.030 ;
        RECT 6.455 30.860 6.955 31.030 ;
        RECT 7.245 30.860 7.745 31.030 ;
        RECT 8.035 30.860 8.535 31.030 ;
        RECT 8.825 30.860 9.325 31.030 ;
        RECT 9.615 30.860 10.115 31.030 ;
        RECT 10.405 30.860 10.905 31.030 ;
        RECT 11.195 30.860 11.695 31.030 ;
        RECT 11.985 30.860 12.485 31.030 ;
        RECT 12.775 30.860 13.275 31.030 ;
        RECT 13.565 30.860 14.065 31.030 ;
        RECT 14.355 30.860 14.855 31.030 ;
        RECT 15.145 30.860 15.645 31.030 ;
        RECT 15.935 30.860 16.435 31.030 ;
        RECT 16.725 30.860 17.225 31.030 ;
        RECT 17.515 30.860 18.015 31.030 ;
        RECT 18.305 30.860 18.805 31.030 ;
        RECT 3.065 29.605 3.235 30.645 ;
        RECT 3.855 29.605 4.025 30.645 ;
        RECT 4.645 29.605 4.815 30.645 ;
        RECT 5.435 29.605 5.605 30.645 ;
        RECT 6.225 29.605 6.395 30.645 ;
        RECT 7.015 29.605 7.185 30.645 ;
        RECT 7.805 29.605 7.975 30.645 ;
        RECT 8.595 29.605 8.765 30.645 ;
        RECT 9.385 29.605 9.555 30.645 ;
        RECT 10.175 29.605 10.345 30.645 ;
        RECT 10.965 29.605 11.135 30.645 ;
        RECT 11.755 29.605 11.925 30.645 ;
        RECT 12.545 29.605 12.715 30.645 ;
        RECT 13.335 29.605 13.505 30.645 ;
        RECT 14.125 29.605 14.295 30.645 ;
        RECT 14.915 29.605 15.085 30.645 ;
        RECT 15.705 29.605 15.875 30.645 ;
        RECT 16.495 29.605 16.665 30.645 ;
        RECT 17.285 29.605 17.455 30.645 ;
        RECT 18.075 29.605 18.245 30.645 ;
        RECT 18.865 29.605 19.035 30.645 ;
        RECT 3.295 29.220 3.795 29.390 ;
        RECT 4.085 29.220 4.585 29.390 ;
        RECT 4.875 29.220 5.375 29.390 ;
        RECT 5.665 29.220 6.165 29.390 ;
        RECT 6.455 29.220 6.955 29.390 ;
        RECT 7.245 29.220 7.745 29.390 ;
        RECT 8.035 29.220 8.535 29.390 ;
        RECT 8.825 29.220 9.325 29.390 ;
        RECT 9.615 29.220 10.115 29.390 ;
        RECT 10.405 29.220 10.905 29.390 ;
        RECT 11.195 29.220 11.695 29.390 ;
        RECT 11.985 29.220 12.485 29.390 ;
        RECT 12.775 29.220 13.275 29.390 ;
        RECT 13.565 29.220 14.065 29.390 ;
        RECT 14.355 29.220 14.855 29.390 ;
        RECT 15.145 29.220 15.645 29.390 ;
        RECT 15.935 29.220 16.435 29.390 ;
        RECT 16.725 29.220 17.225 29.390 ;
        RECT 17.515 29.220 18.015 29.390 ;
        RECT 18.305 29.220 18.805 29.390 ;
        RECT 3.295 28.680 3.795 28.850 ;
        RECT 4.085 28.680 4.585 28.850 ;
        RECT 4.875 28.680 5.375 28.850 ;
        RECT 5.665 28.680 6.165 28.850 ;
        RECT 6.455 28.680 6.955 28.850 ;
        RECT 7.245 28.680 7.745 28.850 ;
        RECT 8.035 28.680 8.535 28.850 ;
        RECT 8.825 28.680 9.325 28.850 ;
        RECT 9.615 28.680 10.115 28.850 ;
        RECT 10.405 28.680 10.905 28.850 ;
        RECT 11.195 28.680 11.695 28.850 ;
        RECT 11.985 28.680 12.485 28.850 ;
        RECT 12.775 28.680 13.275 28.850 ;
        RECT 13.565 28.680 14.065 28.850 ;
        RECT 14.355 28.680 14.855 28.850 ;
        RECT 15.145 28.680 15.645 28.850 ;
        RECT 15.935 28.680 16.435 28.850 ;
        RECT 16.725 28.680 17.225 28.850 ;
        RECT 17.515 28.680 18.015 28.850 ;
        RECT 18.305 28.680 18.805 28.850 ;
        RECT 3.065 27.425 3.235 28.465 ;
        RECT 3.855 27.425 4.025 28.465 ;
        RECT 4.645 27.425 4.815 28.465 ;
        RECT 5.435 27.425 5.605 28.465 ;
        RECT 6.225 27.425 6.395 28.465 ;
        RECT 7.015 27.425 7.185 28.465 ;
        RECT 7.805 27.425 7.975 28.465 ;
        RECT 8.595 27.425 8.765 28.465 ;
        RECT 9.385 27.425 9.555 28.465 ;
        RECT 10.175 27.425 10.345 28.465 ;
        RECT 10.965 27.425 11.135 28.465 ;
        RECT 11.755 27.425 11.925 28.465 ;
        RECT 12.545 27.425 12.715 28.465 ;
        RECT 13.335 27.425 13.505 28.465 ;
        RECT 14.125 27.425 14.295 28.465 ;
        RECT 14.915 27.425 15.085 28.465 ;
        RECT 15.705 27.425 15.875 28.465 ;
        RECT 16.495 27.425 16.665 28.465 ;
        RECT 17.285 27.425 17.455 28.465 ;
        RECT 18.075 27.425 18.245 28.465 ;
        RECT 18.865 27.425 19.035 28.465 ;
        RECT 3.295 27.040 3.795 27.210 ;
        RECT 4.085 27.040 4.585 27.210 ;
        RECT 4.875 27.040 5.375 27.210 ;
        RECT 5.665 27.040 6.165 27.210 ;
        RECT 6.455 27.040 6.955 27.210 ;
        RECT 7.245 27.040 7.745 27.210 ;
        RECT 8.035 27.040 8.535 27.210 ;
        RECT 8.825 27.040 9.325 27.210 ;
        RECT 9.615 27.040 10.115 27.210 ;
        RECT 10.405 27.040 10.905 27.210 ;
        RECT 11.195 27.040 11.695 27.210 ;
        RECT 11.985 27.040 12.485 27.210 ;
        RECT 12.775 27.040 13.275 27.210 ;
        RECT 13.565 27.040 14.065 27.210 ;
        RECT 14.355 27.040 14.855 27.210 ;
        RECT 15.145 27.040 15.645 27.210 ;
        RECT 15.935 27.040 16.435 27.210 ;
        RECT 16.725 27.040 17.225 27.210 ;
        RECT 17.515 27.040 18.015 27.210 ;
        RECT 18.305 27.040 18.805 27.210 ;
        RECT 3.295 26.500 3.795 26.670 ;
        RECT 4.085 26.500 4.585 26.670 ;
        RECT 4.875 26.500 5.375 26.670 ;
        RECT 5.665 26.500 6.165 26.670 ;
        RECT 6.455 26.500 6.955 26.670 ;
        RECT 7.245 26.500 7.745 26.670 ;
        RECT 8.035 26.500 8.535 26.670 ;
        RECT 8.825 26.500 9.325 26.670 ;
        RECT 9.615 26.500 10.115 26.670 ;
        RECT 10.405 26.500 10.905 26.670 ;
        RECT 11.195 26.500 11.695 26.670 ;
        RECT 11.985 26.500 12.485 26.670 ;
        RECT 12.775 26.500 13.275 26.670 ;
        RECT 13.565 26.500 14.065 26.670 ;
        RECT 14.355 26.500 14.855 26.670 ;
        RECT 15.145 26.500 15.645 26.670 ;
        RECT 15.935 26.500 16.435 26.670 ;
        RECT 16.725 26.500 17.225 26.670 ;
        RECT 17.515 26.500 18.015 26.670 ;
        RECT 18.305 26.500 18.805 26.670 ;
        RECT 3.065 25.245 3.235 26.285 ;
        RECT 3.855 25.245 4.025 26.285 ;
        RECT 4.645 25.245 4.815 26.285 ;
        RECT 5.435 25.245 5.605 26.285 ;
        RECT 6.225 25.245 6.395 26.285 ;
        RECT 7.015 25.245 7.185 26.285 ;
        RECT 7.805 25.245 7.975 26.285 ;
        RECT 8.595 25.245 8.765 26.285 ;
        RECT 9.385 25.245 9.555 26.285 ;
        RECT 10.175 25.245 10.345 26.285 ;
        RECT 10.965 25.245 11.135 26.285 ;
        RECT 11.755 25.245 11.925 26.285 ;
        RECT 12.545 25.245 12.715 26.285 ;
        RECT 13.335 25.245 13.505 26.285 ;
        RECT 14.125 25.245 14.295 26.285 ;
        RECT 14.915 25.245 15.085 26.285 ;
        RECT 15.705 25.245 15.875 26.285 ;
        RECT 16.495 25.245 16.665 26.285 ;
        RECT 17.285 25.245 17.455 26.285 ;
        RECT 18.075 25.245 18.245 26.285 ;
        RECT 18.865 25.245 19.035 26.285 ;
        RECT 3.295 24.860 3.795 25.030 ;
        RECT 4.085 24.860 4.585 25.030 ;
        RECT 4.875 24.860 5.375 25.030 ;
        RECT 5.665 24.860 6.165 25.030 ;
        RECT 6.455 24.860 6.955 25.030 ;
        RECT 7.245 24.860 7.745 25.030 ;
        RECT 8.035 24.860 8.535 25.030 ;
        RECT 8.825 24.860 9.325 25.030 ;
        RECT 9.615 24.860 10.115 25.030 ;
        RECT 10.405 24.860 10.905 25.030 ;
        RECT 11.195 24.860 11.695 25.030 ;
        RECT 11.985 24.860 12.485 25.030 ;
        RECT 12.775 24.860 13.275 25.030 ;
        RECT 13.565 24.860 14.065 25.030 ;
        RECT 14.355 24.860 14.855 25.030 ;
        RECT 15.145 24.860 15.645 25.030 ;
        RECT 15.935 24.860 16.435 25.030 ;
        RECT 16.725 24.860 17.225 25.030 ;
        RECT 17.515 24.860 18.015 25.030 ;
        RECT 18.305 24.860 18.805 25.030 ;
        RECT 3.295 24.320 3.795 24.490 ;
        RECT 4.085 24.320 4.585 24.490 ;
        RECT 4.875 24.320 5.375 24.490 ;
        RECT 5.665 24.320 6.165 24.490 ;
        RECT 6.455 24.320 6.955 24.490 ;
        RECT 7.245 24.320 7.745 24.490 ;
        RECT 8.035 24.320 8.535 24.490 ;
        RECT 8.825 24.320 9.325 24.490 ;
        RECT 9.615 24.320 10.115 24.490 ;
        RECT 10.405 24.320 10.905 24.490 ;
        RECT 11.195 24.320 11.695 24.490 ;
        RECT 11.985 24.320 12.485 24.490 ;
        RECT 12.775 24.320 13.275 24.490 ;
        RECT 13.565 24.320 14.065 24.490 ;
        RECT 14.355 24.320 14.855 24.490 ;
        RECT 15.145 24.320 15.645 24.490 ;
        RECT 15.935 24.320 16.435 24.490 ;
        RECT 16.725 24.320 17.225 24.490 ;
        RECT 17.515 24.320 18.015 24.490 ;
        RECT 18.305 24.320 18.805 24.490 ;
        RECT 3.065 23.065 3.235 24.105 ;
        RECT 3.855 23.065 4.025 24.105 ;
        RECT 4.645 23.065 4.815 24.105 ;
        RECT 5.435 23.065 5.605 24.105 ;
        RECT 6.225 23.065 6.395 24.105 ;
        RECT 7.015 23.065 7.185 24.105 ;
        RECT 7.805 23.065 7.975 24.105 ;
        RECT 8.595 23.065 8.765 24.105 ;
        RECT 9.385 23.065 9.555 24.105 ;
        RECT 10.175 23.065 10.345 24.105 ;
        RECT 10.965 23.065 11.135 24.105 ;
        RECT 11.755 23.065 11.925 24.105 ;
        RECT 12.545 23.065 12.715 24.105 ;
        RECT 13.335 23.065 13.505 24.105 ;
        RECT 14.125 23.065 14.295 24.105 ;
        RECT 14.915 23.065 15.085 24.105 ;
        RECT 15.705 23.065 15.875 24.105 ;
        RECT 16.495 23.065 16.665 24.105 ;
        RECT 17.285 23.065 17.455 24.105 ;
        RECT 18.075 23.065 18.245 24.105 ;
        RECT 18.865 23.065 19.035 24.105 ;
        RECT 3.295 22.680 3.795 22.850 ;
        RECT 4.085 22.680 4.585 22.850 ;
        RECT 4.875 22.680 5.375 22.850 ;
        RECT 5.665 22.680 6.165 22.850 ;
        RECT 6.455 22.680 6.955 22.850 ;
        RECT 7.245 22.680 7.745 22.850 ;
        RECT 8.035 22.680 8.535 22.850 ;
        RECT 8.825 22.680 9.325 22.850 ;
        RECT 9.615 22.680 10.115 22.850 ;
        RECT 10.405 22.680 10.905 22.850 ;
        RECT 11.195 22.680 11.695 22.850 ;
        RECT 11.985 22.680 12.485 22.850 ;
        RECT 12.775 22.680 13.275 22.850 ;
        RECT 13.565 22.680 14.065 22.850 ;
        RECT 14.355 22.680 14.855 22.850 ;
        RECT 15.145 22.680 15.645 22.850 ;
        RECT 15.935 22.680 16.435 22.850 ;
        RECT 16.725 22.680 17.225 22.850 ;
        RECT 17.515 22.680 18.015 22.850 ;
        RECT 18.305 22.680 18.805 22.850 ;
        RECT 19.420 22.360 19.865 53.215 ;
        RECT 1.860 21.855 19.865 22.360 ;
        RECT 1.860 19.285 2.710 21.855 ;
        RECT 3.295 21.300 3.795 21.470 ;
        RECT 4.085 21.300 4.585 21.470 ;
        RECT 4.875 21.300 5.375 21.470 ;
        RECT 5.665 21.300 6.165 21.470 ;
        RECT 6.455 21.300 6.955 21.470 ;
        RECT 7.245 21.300 7.745 21.470 ;
        RECT 8.035 21.300 8.535 21.470 ;
        RECT 8.825 21.300 9.325 21.470 ;
        RECT 9.615 21.300 10.115 21.470 ;
        RECT 10.405 21.300 10.905 21.470 ;
        RECT 11.195 21.300 11.695 21.470 ;
        RECT 11.985 21.300 12.485 21.470 ;
        RECT 12.775 21.300 13.275 21.470 ;
        RECT 13.565 21.300 14.065 21.470 ;
        RECT 14.355 21.300 14.855 21.470 ;
        RECT 15.145 21.300 15.645 21.470 ;
        RECT 15.935 21.300 16.435 21.470 ;
        RECT 16.725 21.300 17.225 21.470 ;
        RECT 17.515 21.300 18.015 21.470 ;
        RECT 18.305 21.300 18.805 21.470 ;
        RECT 3.065 20.045 3.235 21.085 ;
        RECT 3.855 20.045 4.025 21.085 ;
        RECT 4.645 20.045 4.815 21.085 ;
        RECT 5.435 20.045 5.605 21.085 ;
        RECT 6.225 20.045 6.395 21.085 ;
        RECT 7.015 20.045 7.185 21.085 ;
        RECT 7.805 20.045 7.975 21.085 ;
        RECT 8.595 20.045 8.765 21.085 ;
        RECT 9.385 20.045 9.555 21.085 ;
        RECT 10.175 20.045 10.345 21.085 ;
        RECT 10.965 20.045 11.135 21.085 ;
        RECT 11.755 20.045 11.925 21.085 ;
        RECT 12.545 20.045 12.715 21.085 ;
        RECT 13.335 20.045 13.505 21.085 ;
        RECT 14.125 20.045 14.295 21.085 ;
        RECT 14.915 20.045 15.085 21.085 ;
        RECT 15.705 20.045 15.875 21.085 ;
        RECT 16.495 20.045 16.665 21.085 ;
        RECT 17.285 20.045 17.455 21.085 ;
        RECT 18.075 20.045 18.245 21.085 ;
        RECT 18.865 20.045 19.035 21.085 ;
        RECT 3.295 19.660 3.795 19.830 ;
        RECT 4.085 19.660 4.585 19.830 ;
        RECT 4.875 19.660 5.375 19.830 ;
        RECT 5.665 19.660 6.165 19.830 ;
        RECT 6.455 19.660 6.955 19.830 ;
        RECT 7.245 19.660 7.745 19.830 ;
        RECT 8.035 19.660 8.535 19.830 ;
        RECT 8.825 19.660 9.325 19.830 ;
        RECT 9.615 19.660 10.115 19.830 ;
        RECT 10.405 19.660 10.905 19.830 ;
        RECT 11.195 19.660 11.695 19.830 ;
        RECT 11.985 19.660 12.485 19.830 ;
        RECT 12.775 19.660 13.275 19.830 ;
        RECT 13.565 19.660 14.065 19.830 ;
        RECT 14.355 19.660 14.855 19.830 ;
        RECT 15.145 19.660 15.645 19.830 ;
        RECT 15.935 19.660 16.435 19.830 ;
        RECT 16.725 19.660 17.225 19.830 ;
        RECT 17.515 19.660 18.015 19.830 ;
        RECT 18.305 19.660 18.805 19.830 ;
        RECT 19.420 19.285 19.865 21.855 ;
        RECT 1.860 18.840 19.865 19.285 ;
        RECT 19.650 18.480 19.845 18.840 ;
        RECT 2.135 18.475 19.895 18.480 ;
        RECT 2.135 17.925 19.955 18.475 ;
        RECT 2.240 15.450 2.795 17.925 ;
        RECT 3.270 17.395 3.770 17.565 ;
        RECT 4.060 17.395 4.560 17.565 ;
        RECT 4.850 17.395 5.350 17.565 ;
        RECT 3.040 16.140 3.210 17.180 ;
        RECT 3.830 16.140 4.000 17.180 ;
        RECT 4.620 16.140 4.790 17.180 ;
        RECT 5.410 16.140 5.580 17.180 ;
        RECT 3.270 15.755 3.770 15.925 ;
        RECT 4.060 15.755 4.560 15.925 ;
        RECT 4.850 15.755 5.350 15.925 ;
        RECT 6.080 15.450 6.250 17.925 ;
        RECT 6.980 17.395 7.480 17.565 ;
        RECT 7.770 17.395 8.270 17.565 ;
        RECT 8.560 17.395 9.060 17.565 ;
        RECT 9.350 17.395 9.850 17.565 ;
        RECT 6.750 16.140 6.920 17.180 ;
        RECT 7.540 16.140 7.710 17.180 ;
        RECT 8.330 16.140 8.500 17.180 ;
        RECT 9.120 16.140 9.290 17.180 ;
        RECT 9.910 16.140 10.080 17.180 ;
        RECT 6.980 15.755 7.480 15.925 ;
        RECT 7.770 15.755 8.270 15.925 ;
        RECT 8.560 15.755 9.060 15.925 ;
        RECT 9.350 15.755 9.850 15.925 ;
        RECT 10.580 15.450 10.750 17.925 ;
        RECT 11.480 17.395 11.980 17.565 ;
        RECT 12.270 17.395 12.770 17.565 ;
        RECT 13.060 17.395 13.560 17.565 ;
        RECT 13.850 17.395 14.350 17.565 ;
        RECT 11.250 16.140 11.420 17.180 ;
        RECT 12.040 16.140 12.210 17.180 ;
        RECT 12.830 16.140 13.000 17.180 ;
        RECT 13.620 16.140 13.790 17.180 ;
        RECT 14.410 16.140 14.580 17.180 ;
        RECT 11.480 15.755 11.980 15.925 ;
        RECT 12.270 15.755 12.770 15.925 ;
        RECT 13.060 15.755 13.560 15.925 ;
        RECT 13.850 15.755 14.350 15.925 ;
        RECT 15.080 15.450 15.250 17.925 ;
        RECT 15.980 17.395 16.480 17.565 ;
        RECT 16.770 17.395 17.270 17.565 ;
        RECT 17.560 17.395 18.060 17.565 ;
        RECT 18.350 17.395 18.850 17.565 ;
        RECT 15.750 16.140 15.920 17.180 ;
        RECT 16.540 16.140 16.710 17.180 ;
        RECT 17.330 16.140 17.500 17.180 ;
        RECT 18.120 16.140 18.290 17.180 ;
        RECT 18.910 16.140 19.080 17.180 ;
        RECT 15.980 15.755 16.480 15.925 ;
        RECT 16.770 15.755 17.270 15.925 ;
        RECT 17.560 15.755 18.060 15.925 ;
        RECT 18.350 15.755 18.850 15.925 ;
        RECT 19.400 15.450 19.955 17.925 ;
        RECT 2.195 14.895 19.955 15.450 ;
        RECT 20.435 15.275 20.940 54.240 ;
        RECT 2.975 13.595 19.525 14.135 ;
        RECT 2.975 11.255 3.515 13.595 ;
        RECT 4.060 13.095 4.560 13.265 ;
        RECT 3.830 11.885 4.000 12.925 ;
        RECT 4.620 11.885 4.790 12.925 ;
        RECT 4.060 11.545 4.560 11.715 ;
        RECT 5.290 11.255 5.480 13.595 ;
        RECT 6.210 13.095 6.710 13.265 ;
        RECT 5.980 11.885 6.150 12.925 ;
        RECT 6.770 11.885 6.940 12.925 ;
        RECT 6.210 11.545 6.710 11.715 ;
        RECT 7.440 11.255 7.630 13.595 ;
        RECT 8.360 13.095 8.860 13.265 ;
        RECT 9.150 13.095 9.650 13.265 ;
        RECT 8.130 11.885 8.300 12.925 ;
        RECT 8.920 11.885 9.090 12.925 ;
        RECT 9.710 11.885 9.880 12.925 ;
        RECT 8.360 11.545 8.860 11.715 ;
        RECT 9.150 11.545 9.650 11.715 ;
        RECT 10.380 11.255 10.570 13.595 ;
        RECT 11.300 13.095 11.800 13.265 ;
        RECT 11.070 11.885 11.240 12.925 ;
        RECT 11.860 11.885 12.030 12.925 ;
        RECT 11.300 11.545 11.800 11.715 ;
        RECT 12.530 11.255 12.720 13.595 ;
        RECT 13.450 13.095 14.350 13.265 ;
        RECT 14.640 13.095 15.540 13.265 ;
        RECT 13.220 11.885 13.390 12.925 ;
        RECT 14.410 11.885 14.580 12.925 ;
        RECT 15.600 11.885 15.770 12.925 ;
        RECT 13.450 11.545 14.350 11.715 ;
        RECT 14.640 11.545 15.540 11.715 ;
        RECT 16.270 11.255 16.460 13.595 ;
        RECT 17.190 13.095 17.690 13.265 ;
        RECT 17.980 13.095 18.480 13.265 ;
        RECT 16.960 11.885 17.130 12.925 ;
        RECT 17.750 11.885 17.920 12.925 ;
        RECT 18.540 11.885 18.710 12.925 ;
        RECT 17.190 11.545 17.690 11.715 ;
        RECT 17.980 11.545 18.480 11.715 ;
        RECT 18.985 11.255 19.525 13.595 ;
        RECT 2.970 10.715 19.525 11.255 ;
        RECT 5.965 10.140 19.525 10.160 ;
        RECT 2.930 9.625 19.525 10.140 ;
        RECT 2.930 8.495 3.435 9.625 ;
        RECT 4.420 9.590 19.525 9.625 ;
        RECT 3.610 8.895 4.100 9.225 ;
        RECT 4.420 8.495 6.075 9.590 ;
        RECT 6.805 9.140 7.305 9.310 ;
        RECT 2.930 8.325 6.075 8.495 ;
        RECT 2.930 7.240 3.435 8.325 ;
        RECT 3.610 7.595 4.100 7.925 ;
        RECT 4.420 7.240 6.075 8.325 ;
        RECT 6.575 7.930 6.745 8.970 ;
        RECT 7.365 7.930 7.535 8.970 ;
        RECT 6.805 7.590 7.305 7.760 ;
        RECT 7.955 7.240 8.465 9.590 ;
        RECT 9.205 9.125 9.705 9.295 ;
        RECT 8.975 7.915 9.145 8.955 ;
        RECT 9.765 7.915 9.935 8.955 ;
        RECT 9.205 7.575 9.705 7.745 ;
        RECT 10.445 7.240 10.955 9.590 ;
        RECT 12.320 8.930 12.730 9.590 ;
        RECT 13.460 9.115 13.960 9.285 ;
        RECT 13.230 8.930 13.400 8.945 ;
        RECT 12.320 7.905 13.400 8.930 ;
        RECT 14.020 7.905 14.190 8.945 ;
        RECT 12.320 7.240 13.270 7.905 ;
        RECT 13.460 7.565 13.960 7.735 ;
        RECT 14.690 7.240 14.880 9.590 ;
        RECT 15.610 9.110 16.110 9.280 ;
        RECT 16.400 9.110 16.900 9.280 ;
        RECT 17.190 9.110 17.690 9.280 ;
        RECT 17.980 9.110 18.480 9.280 ;
        RECT 15.380 7.900 15.550 8.940 ;
        RECT 16.170 7.900 16.340 8.940 ;
        RECT 16.960 7.900 17.130 8.940 ;
        RECT 17.750 7.900 17.920 8.940 ;
        RECT 18.540 7.900 18.710 8.940 ;
        RECT 15.610 7.560 16.110 7.730 ;
        RECT 16.400 7.560 16.900 7.730 ;
        RECT 17.190 7.560 17.690 7.730 ;
        RECT 17.980 7.560 18.480 7.730 ;
        RECT 18.955 7.240 19.525 9.590 ;
        RECT 2.930 6.670 19.525 7.240 ;
        RECT 2.210 5.475 20.075 6.015 ;
        RECT 2.210 -4.740 2.685 5.475 ;
        RECT 3.025 4.680 5.185 5.030 ;
        RECT 16.685 4.680 18.845 5.030 ;
        RECT 3.025 3.850 5.185 4.200 ;
        RECT 16.685 3.850 18.845 4.200 ;
        RECT 3.025 3.020 5.185 3.370 ;
        RECT 16.685 3.020 18.845 3.370 ;
        RECT 3.025 2.190 5.185 2.540 ;
        RECT 16.685 2.190 18.845 2.540 ;
        RECT 3.025 1.360 5.185 1.710 ;
        RECT 16.685 1.360 18.845 1.710 ;
        RECT 3.025 0.530 5.185 0.880 ;
        RECT 16.685 0.530 18.845 0.880 ;
        RECT 3.025 -0.300 5.185 0.050 ;
        RECT 16.685 -0.300 18.845 0.050 ;
        RECT 3.025 -1.130 5.185 -0.780 ;
        RECT 16.685 -1.130 18.845 -0.780 ;
        RECT 3.025 -1.960 5.185 -1.610 ;
        RECT 16.685 -1.960 18.845 -1.610 ;
        RECT 3.025 -2.790 5.185 -2.440 ;
        RECT 16.685 -2.790 18.845 -2.440 ;
        RECT 3.025 -3.620 5.185 -3.270 ;
        RECT 16.685 -3.620 18.845 -3.270 ;
        RECT 3.025 -4.450 5.185 -4.100 ;
        RECT 16.685 -4.450 18.845 -4.100 ;
        RECT 19.325 -4.740 20.075 5.475 ;
        RECT 2.210 -5.270 20.075 -4.740 ;
        RECT 20.670 -6.075 20.840 15.275 ;
        RECT 0.895 -6.635 20.975 -6.075 ;
        RECT 21.390 -6.970 21.885 55.145 ;
        RECT 0.000 -7.480 21.885 -6.970 ;
      LAYER met1 ;
        RECT 0.000 55.145 21.885 55.645 ;
        RECT 0.000 -6.735 0.540 55.145 ;
        RECT 0.895 54.695 1.415 54.715 ;
        RECT 0.895 54.240 20.940 54.695 ;
        RECT 0.895 22.465 1.415 54.240 ;
        RECT 1.765 53.665 2.290 54.240 ;
        RECT 19.535 53.670 20.060 54.240 ;
        RECT 19.535 53.665 20.070 53.670 ;
        RECT 1.765 53.660 20.070 53.665 ;
        RECT 1.750 53.220 20.070 53.660 ;
        RECT 1.750 22.465 2.285 53.220 ;
        RECT 0.895 21.875 2.285 22.465 ;
        RECT 0.895 18.465 1.415 21.875 ;
        RECT 1.750 18.465 2.285 21.875 ;
        RECT 2.525 52.840 3.775 52.860 ;
        RECT 4.105 52.840 4.565 52.860 ;
        RECT 4.895 52.840 5.355 52.860 ;
        RECT 5.685 52.840 6.145 52.860 ;
        RECT 6.475 52.840 6.935 52.860 ;
        RECT 7.265 52.840 7.725 52.860 ;
        RECT 8.055 52.840 8.515 52.860 ;
        RECT 8.845 52.840 9.305 52.860 ;
        RECT 9.635 52.840 10.095 52.860 ;
        RECT 10.425 52.840 10.885 52.860 ;
        RECT 11.215 52.840 11.675 52.860 ;
        RECT 12.005 52.840 12.465 52.860 ;
        RECT 12.795 52.840 13.255 52.860 ;
        RECT 13.585 52.840 14.045 52.860 ;
        RECT 14.375 52.840 14.835 52.860 ;
        RECT 15.165 52.840 15.625 52.860 ;
        RECT 15.955 52.840 16.415 52.860 ;
        RECT 16.745 52.840 17.205 52.860 ;
        RECT 17.535 52.840 17.995 52.860 ;
        RECT 18.325 52.840 18.785 52.860 ;
        RECT 2.525 52.655 18.825 52.840 ;
        RECT 2.525 52.630 3.775 52.655 ;
        RECT 4.105 52.630 4.565 52.655 ;
        RECT 4.895 52.630 5.355 52.655 ;
        RECT 5.685 52.630 6.145 52.655 ;
        RECT 6.475 52.630 6.935 52.655 ;
        RECT 7.265 52.630 7.725 52.655 ;
        RECT 8.055 52.630 8.515 52.655 ;
        RECT 8.845 52.630 9.305 52.655 ;
        RECT 9.635 52.630 10.095 52.655 ;
        RECT 10.425 52.630 10.885 52.655 ;
        RECT 11.215 52.630 11.675 52.655 ;
        RECT 12.005 52.630 12.465 52.655 ;
        RECT 12.795 52.630 13.255 52.655 ;
        RECT 13.585 52.630 14.045 52.655 ;
        RECT 14.375 52.630 14.835 52.655 ;
        RECT 15.165 52.630 15.625 52.655 ;
        RECT 15.955 52.630 16.415 52.655 ;
        RECT 16.745 52.630 17.205 52.655 ;
        RECT 17.535 52.630 17.995 52.655 ;
        RECT 18.325 52.630 18.785 52.655 ;
        RECT 2.525 51.220 2.760 52.630 ;
        RECT 3.020 51.815 3.280 52.485 ;
        RECT 3.035 51.425 3.265 51.815 ;
        RECT 3.460 51.220 3.620 52.630 ;
        RECT 3.825 52.045 4.055 52.425 ;
        RECT 3.810 51.375 4.070 52.045 ;
        RECT 4.250 51.220 4.410 52.630 ;
        RECT 4.600 51.815 4.860 52.485 ;
        RECT 4.615 51.425 4.845 51.815 ;
        RECT 5.040 51.220 5.200 52.630 ;
        RECT 5.405 52.045 5.635 52.425 ;
        RECT 5.390 51.375 5.650 52.045 ;
        RECT 5.830 51.220 5.990 52.630 ;
        RECT 6.180 51.815 6.440 52.485 ;
        RECT 6.195 51.425 6.425 51.815 ;
        RECT 6.620 51.220 6.780 52.630 ;
        RECT 6.985 52.045 7.215 52.425 ;
        RECT 6.970 51.375 7.230 52.045 ;
        RECT 7.410 51.220 7.570 52.630 ;
        RECT 7.760 51.815 8.020 52.485 ;
        RECT 7.775 51.425 8.005 51.815 ;
        RECT 8.200 51.220 8.360 52.630 ;
        RECT 8.565 52.045 8.795 52.425 ;
        RECT 8.550 51.375 8.810 52.045 ;
        RECT 8.990 51.220 9.150 52.630 ;
        RECT 9.340 51.815 9.600 52.485 ;
        RECT 9.355 51.425 9.585 51.815 ;
        RECT 9.780 51.220 9.940 52.630 ;
        RECT 10.145 52.045 10.375 52.425 ;
        RECT 10.130 51.375 10.390 52.045 ;
        RECT 10.570 51.220 10.730 52.630 ;
        RECT 10.920 51.815 11.180 52.485 ;
        RECT 10.935 51.425 11.165 51.815 ;
        RECT 11.360 51.220 11.520 52.630 ;
        RECT 11.725 52.045 11.955 52.425 ;
        RECT 11.710 51.375 11.970 52.045 ;
        RECT 12.150 51.220 12.310 52.630 ;
        RECT 12.500 51.815 12.760 52.485 ;
        RECT 12.515 51.425 12.745 51.815 ;
        RECT 12.940 51.220 13.100 52.630 ;
        RECT 13.305 52.045 13.535 52.425 ;
        RECT 13.290 51.375 13.550 52.045 ;
        RECT 13.730 51.220 13.890 52.630 ;
        RECT 14.080 51.815 14.340 52.485 ;
        RECT 14.095 51.425 14.325 51.815 ;
        RECT 14.520 51.220 14.680 52.630 ;
        RECT 14.885 52.045 15.115 52.425 ;
        RECT 14.870 51.375 15.130 52.045 ;
        RECT 15.310 51.220 15.470 52.630 ;
        RECT 15.660 51.815 15.920 52.485 ;
        RECT 15.675 51.425 15.905 51.815 ;
        RECT 16.100 51.220 16.260 52.630 ;
        RECT 16.465 52.045 16.695 52.425 ;
        RECT 16.450 51.375 16.710 52.045 ;
        RECT 16.890 51.220 17.050 52.630 ;
        RECT 17.240 51.815 17.500 52.485 ;
        RECT 17.255 51.425 17.485 51.815 ;
        RECT 17.680 51.220 17.840 52.630 ;
        RECT 18.045 52.045 18.275 52.425 ;
        RECT 18.030 51.375 18.290 52.045 ;
        RECT 18.470 51.220 18.630 52.630 ;
        RECT 18.820 51.815 19.080 52.485 ;
        RECT 18.835 51.425 19.065 51.815 ;
        RECT 2.525 51.200 3.775 51.220 ;
        RECT 4.105 51.200 4.565 51.220 ;
        RECT 4.895 51.200 5.355 51.220 ;
        RECT 5.685 51.200 6.145 51.220 ;
        RECT 6.475 51.200 6.935 51.220 ;
        RECT 7.265 51.200 7.725 51.220 ;
        RECT 8.055 51.200 8.515 51.220 ;
        RECT 8.845 51.200 9.305 51.220 ;
        RECT 9.635 51.200 10.095 51.220 ;
        RECT 10.425 51.200 10.885 51.220 ;
        RECT 11.215 51.200 11.675 51.220 ;
        RECT 12.005 51.200 12.465 51.220 ;
        RECT 12.795 51.200 13.255 51.220 ;
        RECT 13.585 51.200 14.045 51.220 ;
        RECT 14.375 51.200 14.835 51.220 ;
        RECT 15.165 51.200 15.625 51.220 ;
        RECT 15.955 51.200 16.415 51.220 ;
        RECT 16.745 51.200 17.205 51.220 ;
        RECT 17.535 51.200 17.995 51.220 ;
        RECT 18.325 51.200 18.785 51.220 ;
        RECT 2.525 51.015 18.785 51.200 ;
        RECT 2.525 50.990 3.775 51.015 ;
        RECT 4.105 50.990 4.565 51.015 ;
        RECT 4.895 50.990 5.355 51.015 ;
        RECT 5.685 50.990 6.145 51.015 ;
        RECT 6.475 50.990 6.935 51.015 ;
        RECT 7.265 50.990 7.725 51.015 ;
        RECT 8.055 50.990 8.515 51.015 ;
        RECT 8.845 50.990 9.305 51.015 ;
        RECT 9.635 50.990 10.095 51.015 ;
        RECT 10.425 50.990 10.885 51.015 ;
        RECT 11.215 50.990 11.675 51.015 ;
        RECT 12.005 50.990 12.465 51.015 ;
        RECT 12.795 50.990 13.255 51.015 ;
        RECT 13.585 50.990 14.045 51.015 ;
        RECT 14.375 50.990 14.835 51.015 ;
        RECT 15.165 50.990 15.625 51.015 ;
        RECT 15.955 50.990 16.415 51.015 ;
        RECT 16.745 50.990 17.205 51.015 ;
        RECT 17.535 50.990 17.995 51.015 ;
        RECT 18.325 50.990 18.785 51.015 ;
        RECT 2.525 50.680 2.760 50.990 ;
        RECT 3.460 50.680 3.620 50.990 ;
        RECT 4.250 50.680 4.410 50.990 ;
        RECT 5.040 50.680 5.200 50.990 ;
        RECT 5.830 50.680 5.990 50.990 ;
        RECT 6.620 50.680 6.780 50.990 ;
        RECT 7.410 50.680 7.570 50.990 ;
        RECT 8.200 50.680 8.360 50.990 ;
        RECT 8.990 50.680 9.150 50.990 ;
        RECT 9.780 50.680 9.940 50.990 ;
        RECT 10.570 50.680 10.730 50.990 ;
        RECT 11.360 50.680 11.520 50.990 ;
        RECT 12.150 50.680 12.310 50.990 ;
        RECT 12.940 50.680 13.100 50.990 ;
        RECT 13.730 50.680 13.890 50.990 ;
        RECT 14.520 50.680 14.680 50.990 ;
        RECT 15.310 50.680 15.470 50.990 ;
        RECT 16.100 50.680 16.260 50.990 ;
        RECT 16.890 50.680 17.050 50.990 ;
        RECT 17.680 50.680 17.840 50.990 ;
        RECT 18.470 50.680 18.630 50.990 ;
        RECT 2.525 50.660 3.775 50.680 ;
        RECT 4.105 50.660 4.565 50.680 ;
        RECT 4.895 50.660 5.355 50.680 ;
        RECT 5.685 50.660 6.145 50.680 ;
        RECT 6.475 50.660 6.935 50.680 ;
        RECT 7.265 50.660 7.725 50.680 ;
        RECT 8.055 50.660 8.515 50.680 ;
        RECT 8.845 50.660 9.305 50.680 ;
        RECT 9.635 50.660 10.095 50.680 ;
        RECT 10.425 50.660 10.885 50.680 ;
        RECT 11.215 50.660 11.675 50.680 ;
        RECT 12.005 50.660 12.465 50.680 ;
        RECT 12.795 50.660 13.255 50.680 ;
        RECT 13.585 50.660 14.045 50.680 ;
        RECT 14.375 50.660 14.835 50.680 ;
        RECT 15.165 50.660 15.625 50.680 ;
        RECT 15.955 50.660 16.415 50.680 ;
        RECT 16.745 50.660 17.205 50.680 ;
        RECT 17.535 50.660 17.995 50.680 ;
        RECT 18.325 50.660 18.785 50.680 ;
        RECT 2.525 50.475 18.825 50.660 ;
        RECT 2.525 50.450 3.775 50.475 ;
        RECT 4.105 50.450 4.565 50.475 ;
        RECT 4.895 50.450 5.355 50.475 ;
        RECT 5.685 50.450 6.145 50.475 ;
        RECT 6.475 50.450 6.935 50.475 ;
        RECT 7.265 50.450 7.725 50.475 ;
        RECT 8.055 50.450 8.515 50.475 ;
        RECT 8.845 50.450 9.305 50.475 ;
        RECT 9.635 50.450 10.095 50.475 ;
        RECT 10.425 50.450 10.885 50.475 ;
        RECT 11.215 50.450 11.675 50.475 ;
        RECT 12.005 50.450 12.465 50.475 ;
        RECT 12.795 50.450 13.255 50.475 ;
        RECT 13.585 50.450 14.045 50.475 ;
        RECT 14.375 50.450 14.835 50.475 ;
        RECT 15.165 50.450 15.625 50.475 ;
        RECT 15.955 50.450 16.415 50.475 ;
        RECT 16.745 50.450 17.205 50.475 ;
        RECT 17.535 50.450 17.995 50.475 ;
        RECT 18.325 50.450 18.785 50.475 ;
        RECT 2.525 49.040 2.760 50.450 ;
        RECT 3.020 49.635 3.280 50.305 ;
        RECT 3.035 49.245 3.265 49.635 ;
        RECT 3.460 49.040 3.620 50.450 ;
        RECT 3.825 49.865 4.055 50.245 ;
        RECT 3.810 49.195 4.070 49.865 ;
        RECT 4.250 49.040 4.410 50.450 ;
        RECT 4.600 49.635 4.860 50.305 ;
        RECT 4.615 49.245 4.845 49.635 ;
        RECT 5.040 49.040 5.200 50.450 ;
        RECT 5.405 49.865 5.635 50.245 ;
        RECT 5.390 49.195 5.650 49.865 ;
        RECT 5.830 49.040 5.990 50.450 ;
        RECT 6.180 49.635 6.440 50.305 ;
        RECT 6.195 49.245 6.425 49.635 ;
        RECT 6.620 49.040 6.780 50.450 ;
        RECT 6.985 49.865 7.215 50.245 ;
        RECT 6.970 49.195 7.230 49.865 ;
        RECT 7.410 49.040 7.570 50.450 ;
        RECT 7.760 49.635 8.020 50.305 ;
        RECT 7.775 49.245 8.005 49.635 ;
        RECT 8.200 49.040 8.360 50.450 ;
        RECT 8.565 49.865 8.795 50.245 ;
        RECT 8.550 49.195 8.810 49.865 ;
        RECT 8.990 49.040 9.150 50.450 ;
        RECT 9.340 49.635 9.600 50.305 ;
        RECT 9.355 49.245 9.585 49.635 ;
        RECT 9.780 49.040 9.940 50.450 ;
        RECT 10.145 49.865 10.375 50.245 ;
        RECT 10.130 49.195 10.390 49.865 ;
        RECT 10.570 49.040 10.730 50.450 ;
        RECT 10.920 49.635 11.180 50.305 ;
        RECT 10.935 49.245 11.165 49.635 ;
        RECT 11.360 49.040 11.520 50.450 ;
        RECT 11.725 49.865 11.955 50.245 ;
        RECT 11.710 49.195 11.970 49.865 ;
        RECT 12.150 49.040 12.310 50.450 ;
        RECT 12.500 49.635 12.760 50.305 ;
        RECT 12.515 49.245 12.745 49.635 ;
        RECT 12.940 49.040 13.100 50.450 ;
        RECT 13.305 49.865 13.535 50.245 ;
        RECT 13.290 49.195 13.550 49.865 ;
        RECT 13.730 49.040 13.890 50.450 ;
        RECT 14.080 49.635 14.340 50.305 ;
        RECT 14.095 49.245 14.325 49.635 ;
        RECT 14.520 49.040 14.680 50.450 ;
        RECT 14.885 49.865 15.115 50.245 ;
        RECT 14.870 49.195 15.130 49.865 ;
        RECT 15.310 49.040 15.470 50.450 ;
        RECT 15.660 49.635 15.920 50.305 ;
        RECT 15.675 49.245 15.905 49.635 ;
        RECT 16.100 49.040 16.260 50.450 ;
        RECT 16.465 49.865 16.695 50.245 ;
        RECT 16.450 49.195 16.710 49.865 ;
        RECT 16.890 49.040 17.050 50.450 ;
        RECT 17.240 49.635 17.500 50.305 ;
        RECT 17.255 49.245 17.485 49.635 ;
        RECT 17.680 49.040 17.840 50.450 ;
        RECT 18.045 49.865 18.275 50.245 ;
        RECT 18.030 49.195 18.290 49.865 ;
        RECT 18.470 49.040 18.630 50.450 ;
        RECT 18.820 49.635 19.080 50.305 ;
        RECT 18.835 49.245 19.065 49.635 ;
        RECT 2.525 49.020 3.775 49.040 ;
        RECT 4.105 49.020 4.565 49.040 ;
        RECT 4.895 49.020 5.355 49.040 ;
        RECT 5.685 49.020 6.145 49.040 ;
        RECT 6.475 49.020 6.935 49.040 ;
        RECT 7.265 49.020 7.725 49.040 ;
        RECT 8.055 49.020 8.515 49.040 ;
        RECT 8.845 49.020 9.305 49.040 ;
        RECT 9.635 49.020 10.095 49.040 ;
        RECT 10.425 49.020 10.885 49.040 ;
        RECT 11.215 49.020 11.675 49.040 ;
        RECT 12.005 49.020 12.465 49.040 ;
        RECT 12.795 49.020 13.255 49.040 ;
        RECT 13.585 49.020 14.045 49.040 ;
        RECT 14.375 49.020 14.835 49.040 ;
        RECT 15.165 49.020 15.625 49.040 ;
        RECT 15.955 49.020 16.415 49.040 ;
        RECT 16.745 49.020 17.205 49.040 ;
        RECT 17.535 49.020 17.995 49.040 ;
        RECT 18.325 49.020 18.785 49.040 ;
        RECT 2.525 48.835 18.785 49.020 ;
        RECT 2.525 48.810 3.775 48.835 ;
        RECT 4.105 48.810 4.565 48.835 ;
        RECT 4.895 48.810 5.355 48.835 ;
        RECT 5.685 48.810 6.145 48.835 ;
        RECT 6.475 48.810 6.935 48.835 ;
        RECT 7.265 48.810 7.725 48.835 ;
        RECT 8.055 48.810 8.515 48.835 ;
        RECT 8.845 48.810 9.305 48.835 ;
        RECT 9.635 48.810 10.095 48.835 ;
        RECT 10.425 48.810 10.885 48.835 ;
        RECT 11.215 48.810 11.675 48.835 ;
        RECT 12.005 48.810 12.465 48.835 ;
        RECT 12.795 48.810 13.255 48.835 ;
        RECT 13.585 48.810 14.045 48.835 ;
        RECT 14.375 48.810 14.835 48.835 ;
        RECT 15.165 48.810 15.625 48.835 ;
        RECT 15.955 48.810 16.415 48.835 ;
        RECT 16.745 48.810 17.205 48.835 ;
        RECT 17.535 48.810 17.995 48.835 ;
        RECT 18.325 48.810 18.785 48.835 ;
        RECT 2.525 48.500 2.760 48.810 ;
        RECT 3.460 48.500 3.620 48.810 ;
        RECT 4.250 48.500 4.410 48.810 ;
        RECT 5.040 48.500 5.200 48.810 ;
        RECT 5.830 48.500 5.990 48.810 ;
        RECT 6.620 48.500 6.780 48.810 ;
        RECT 7.410 48.500 7.570 48.810 ;
        RECT 8.200 48.500 8.360 48.810 ;
        RECT 8.990 48.500 9.150 48.810 ;
        RECT 9.780 48.500 9.940 48.810 ;
        RECT 10.570 48.500 10.730 48.810 ;
        RECT 11.360 48.500 11.520 48.810 ;
        RECT 12.150 48.500 12.310 48.810 ;
        RECT 12.940 48.500 13.100 48.810 ;
        RECT 13.730 48.500 13.890 48.810 ;
        RECT 14.520 48.500 14.680 48.810 ;
        RECT 15.310 48.500 15.470 48.810 ;
        RECT 16.100 48.500 16.260 48.810 ;
        RECT 16.890 48.500 17.050 48.810 ;
        RECT 17.680 48.500 17.840 48.810 ;
        RECT 18.470 48.500 18.630 48.810 ;
        RECT 2.525 48.480 3.775 48.500 ;
        RECT 4.105 48.480 4.565 48.500 ;
        RECT 4.895 48.480 5.355 48.500 ;
        RECT 5.685 48.480 6.145 48.500 ;
        RECT 6.475 48.480 6.935 48.500 ;
        RECT 7.265 48.480 7.725 48.500 ;
        RECT 8.055 48.480 8.515 48.500 ;
        RECT 8.845 48.480 9.305 48.500 ;
        RECT 9.635 48.480 10.095 48.500 ;
        RECT 10.425 48.480 10.885 48.500 ;
        RECT 11.215 48.480 11.675 48.500 ;
        RECT 12.005 48.480 12.465 48.500 ;
        RECT 12.795 48.480 13.255 48.500 ;
        RECT 13.585 48.480 14.045 48.500 ;
        RECT 14.375 48.480 14.835 48.500 ;
        RECT 15.165 48.480 15.625 48.500 ;
        RECT 15.955 48.480 16.415 48.500 ;
        RECT 16.745 48.480 17.205 48.500 ;
        RECT 17.535 48.480 17.995 48.500 ;
        RECT 18.325 48.480 18.785 48.500 ;
        RECT 2.525 48.295 18.825 48.480 ;
        RECT 2.525 48.270 3.775 48.295 ;
        RECT 4.105 48.270 4.565 48.295 ;
        RECT 4.895 48.270 5.355 48.295 ;
        RECT 5.685 48.270 6.145 48.295 ;
        RECT 6.475 48.270 6.935 48.295 ;
        RECT 7.265 48.270 7.725 48.295 ;
        RECT 8.055 48.270 8.515 48.295 ;
        RECT 8.845 48.270 9.305 48.295 ;
        RECT 9.635 48.270 10.095 48.295 ;
        RECT 10.425 48.270 10.885 48.295 ;
        RECT 11.215 48.270 11.675 48.295 ;
        RECT 12.005 48.270 12.465 48.295 ;
        RECT 12.795 48.270 13.255 48.295 ;
        RECT 13.585 48.270 14.045 48.295 ;
        RECT 14.375 48.270 14.835 48.295 ;
        RECT 15.165 48.270 15.625 48.295 ;
        RECT 15.955 48.270 16.415 48.295 ;
        RECT 16.745 48.270 17.205 48.295 ;
        RECT 17.535 48.270 17.995 48.295 ;
        RECT 18.325 48.270 18.785 48.295 ;
        RECT 2.525 46.860 2.760 48.270 ;
        RECT 3.020 47.455 3.280 48.125 ;
        RECT 3.035 47.065 3.265 47.455 ;
        RECT 3.460 46.860 3.620 48.270 ;
        RECT 3.825 47.685 4.055 48.065 ;
        RECT 3.810 47.015 4.070 47.685 ;
        RECT 4.250 46.860 4.410 48.270 ;
        RECT 4.600 47.455 4.860 48.125 ;
        RECT 4.615 47.065 4.845 47.455 ;
        RECT 5.040 46.860 5.200 48.270 ;
        RECT 5.405 47.685 5.635 48.065 ;
        RECT 5.390 47.015 5.650 47.685 ;
        RECT 5.830 46.860 5.990 48.270 ;
        RECT 6.180 47.455 6.440 48.125 ;
        RECT 6.195 47.065 6.425 47.455 ;
        RECT 6.620 46.860 6.780 48.270 ;
        RECT 6.985 47.685 7.215 48.065 ;
        RECT 6.970 47.015 7.230 47.685 ;
        RECT 7.410 46.860 7.570 48.270 ;
        RECT 7.760 47.455 8.020 48.125 ;
        RECT 7.775 47.065 8.005 47.455 ;
        RECT 8.200 46.860 8.360 48.270 ;
        RECT 8.565 47.685 8.795 48.065 ;
        RECT 8.550 47.015 8.810 47.685 ;
        RECT 8.990 46.860 9.150 48.270 ;
        RECT 9.340 47.455 9.600 48.125 ;
        RECT 9.355 47.065 9.585 47.455 ;
        RECT 9.780 46.860 9.940 48.270 ;
        RECT 10.145 47.685 10.375 48.065 ;
        RECT 10.130 47.015 10.390 47.685 ;
        RECT 10.570 46.860 10.730 48.270 ;
        RECT 10.920 47.455 11.180 48.125 ;
        RECT 10.935 47.065 11.165 47.455 ;
        RECT 11.360 46.860 11.520 48.270 ;
        RECT 11.725 47.685 11.955 48.065 ;
        RECT 11.710 47.015 11.970 47.685 ;
        RECT 12.150 46.860 12.310 48.270 ;
        RECT 12.500 47.455 12.760 48.125 ;
        RECT 12.515 47.065 12.745 47.455 ;
        RECT 12.940 46.860 13.100 48.270 ;
        RECT 13.305 47.685 13.535 48.065 ;
        RECT 13.290 47.015 13.550 47.685 ;
        RECT 13.730 46.860 13.890 48.270 ;
        RECT 14.080 47.455 14.340 48.125 ;
        RECT 14.095 47.065 14.325 47.455 ;
        RECT 14.520 46.860 14.680 48.270 ;
        RECT 14.885 47.685 15.115 48.065 ;
        RECT 14.870 47.015 15.130 47.685 ;
        RECT 15.310 46.860 15.470 48.270 ;
        RECT 15.660 47.455 15.920 48.125 ;
        RECT 15.675 47.065 15.905 47.455 ;
        RECT 16.100 46.860 16.260 48.270 ;
        RECT 16.465 47.685 16.695 48.065 ;
        RECT 16.450 47.015 16.710 47.685 ;
        RECT 16.890 46.860 17.050 48.270 ;
        RECT 17.240 47.455 17.500 48.125 ;
        RECT 17.255 47.065 17.485 47.455 ;
        RECT 17.680 46.860 17.840 48.270 ;
        RECT 18.045 47.685 18.275 48.065 ;
        RECT 18.030 47.015 18.290 47.685 ;
        RECT 18.470 46.860 18.630 48.270 ;
        RECT 18.820 47.455 19.080 48.125 ;
        RECT 18.835 47.065 19.065 47.455 ;
        RECT 2.525 46.840 3.775 46.860 ;
        RECT 4.105 46.840 4.565 46.860 ;
        RECT 4.895 46.840 5.355 46.860 ;
        RECT 5.685 46.840 6.145 46.860 ;
        RECT 6.475 46.840 6.935 46.860 ;
        RECT 7.265 46.840 7.725 46.860 ;
        RECT 8.055 46.840 8.515 46.860 ;
        RECT 8.845 46.840 9.305 46.860 ;
        RECT 9.635 46.840 10.095 46.860 ;
        RECT 10.425 46.840 10.885 46.860 ;
        RECT 11.215 46.840 11.675 46.860 ;
        RECT 12.005 46.840 12.465 46.860 ;
        RECT 12.795 46.840 13.255 46.860 ;
        RECT 13.585 46.840 14.045 46.860 ;
        RECT 14.375 46.840 14.835 46.860 ;
        RECT 15.165 46.840 15.625 46.860 ;
        RECT 15.955 46.840 16.415 46.860 ;
        RECT 16.745 46.840 17.205 46.860 ;
        RECT 17.535 46.840 17.995 46.860 ;
        RECT 18.325 46.840 18.785 46.860 ;
        RECT 2.525 46.655 18.785 46.840 ;
        RECT 2.525 46.630 3.775 46.655 ;
        RECT 4.105 46.630 4.565 46.655 ;
        RECT 4.895 46.630 5.355 46.655 ;
        RECT 5.685 46.630 6.145 46.655 ;
        RECT 6.475 46.630 6.935 46.655 ;
        RECT 7.265 46.630 7.725 46.655 ;
        RECT 8.055 46.630 8.515 46.655 ;
        RECT 8.845 46.630 9.305 46.655 ;
        RECT 9.635 46.630 10.095 46.655 ;
        RECT 10.425 46.630 10.885 46.655 ;
        RECT 11.215 46.630 11.675 46.655 ;
        RECT 12.005 46.630 12.465 46.655 ;
        RECT 12.795 46.630 13.255 46.655 ;
        RECT 13.585 46.630 14.045 46.655 ;
        RECT 14.375 46.630 14.835 46.655 ;
        RECT 15.165 46.630 15.625 46.655 ;
        RECT 15.955 46.630 16.415 46.655 ;
        RECT 16.745 46.630 17.205 46.655 ;
        RECT 17.535 46.630 17.995 46.655 ;
        RECT 18.325 46.630 18.785 46.655 ;
        RECT 2.525 46.320 2.760 46.630 ;
        RECT 3.460 46.320 3.620 46.630 ;
        RECT 4.250 46.320 4.410 46.630 ;
        RECT 5.040 46.320 5.200 46.630 ;
        RECT 5.830 46.320 5.990 46.630 ;
        RECT 6.620 46.320 6.780 46.630 ;
        RECT 7.410 46.320 7.570 46.630 ;
        RECT 8.200 46.320 8.360 46.630 ;
        RECT 8.990 46.320 9.150 46.630 ;
        RECT 9.780 46.320 9.940 46.630 ;
        RECT 10.570 46.320 10.730 46.630 ;
        RECT 11.360 46.320 11.520 46.630 ;
        RECT 12.150 46.320 12.310 46.630 ;
        RECT 12.940 46.320 13.100 46.630 ;
        RECT 13.730 46.320 13.890 46.630 ;
        RECT 14.520 46.320 14.680 46.630 ;
        RECT 15.310 46.320 15.470 46.630 ;
        RECT 16.100 46.320 16.260 46.630 ;
        RECT 16.890 46.320 17.050 46.630 ;
        RECT 17.680 46.320 17.840 46.630 ;
        RECT 18.470 46.320 18.630 46.630 ;
        RECT 2.525 46.300 3.775 46.320 ;
        RECT 4.105 46.300 4.565 46.320 ;
        RECT 4.895 46.300 5.355 46.320 ;
        RECT 5.685 46.300 6.145 46.320 ;
        RECT 6.475 46.300 6.935 46.320 ;
        RECT 7.265 46.300 7.725 46.320 ;
        RECT 8.055 46.300 8.515 46.320 ;
        RECT 8.845 46.300 9.305 46.320 ;
        RECT 9.635 46.300 10.095 46.320 ;
        RECT 10.425 46.300 10.885 46.320 ;
        RECT 11.215 46.300 11.675 46.320 ;
        RECT 12.005 46.300 12.465 46.320 ;
        RECT 12.795 46.300 13.255 46.320 ;
        RECT 13.585 46.300 14.045 46.320 ;
        RECT 14.375 46.300 14.835 46.320 ;
        RECT 15.165 46.300 15.625 46.320 ;
        RECT 15.955 46.300 16.415 46.320 ;
        RECT 16.745 46.300 17.205 46.320 ;
        RECT 17.535 46.300 17.995 46.320 ;
        RECT 18.325 46.300 18.785 46.320 ;
        RECT 2.525 46.115 18.825 46.300 ;
        RECT 2.525 46.090 3.775 46.115 ;
        RECT 4.105 46.090 4.565 46.115 ;
        RECT 4.895 46.090 5.355 46.115 ;
        RECT 5.685 46.090 6.145 46.115 ;
        RECT 6.475 46.090 6.935 46.115 ;
        RECT 7.265 46.090 7.725 46.115 ;
        RECT 8.055 46.090 8.515 46.115 ;
        RECT 8.845 46.090 9.305 46.115 ;
        RECT 9.635 46.090 10.095 46.115 ;
        RECT 10.425 46.090 10.885 46.115 ;
        RECT 11.215 46.090 11.675 46.115 ;
        RECT 12.005 46.090 12.465 46.115 ;
        RECT 12.795 46.090 13.255 46.115 ;
        RECT 13.585 46.090 14.045 46.115 ;
        RECT 14.375 46.090 14.835 46.115 ;
        RECT 15.165 46.090 15.625 46.115 ;
        RECT 15.955 46.090 16.415 46.115 ;
        RECT 16.745 46.090 17.205 46.115 ;
        RECT 17.535 46.090 17.995 46.115 ;
        RECT 18.325 46.090 18.785 46.115 ;
        RECT 2.525 44.680 2.760 46.090 ;
        RECT 3.020 45.275 3.280 45.945 ;
        RECT 3.035 44.885 3.265 45.275 ;
        RECT 3.460 44.680 3.620 46.090 ;
        RECT 3.825 45.505 4.055 45.885 ;
        RECT 3.810 44.835 4.070 45.505 ;
        RECT 4.250 44.680 4.410 46.090 ;
        RECT 4.600 45.275 4.860 45.945 ;
        RECT 4.615 44.885 4.845 45.275 ;
        RECT 5.040 44.680 5.200 46.090 ;
        RECT 5.405 45.505 5.635 45.885 ;
        RECT 5.390 44.835 5.650 45.505 ;
        RECT 5.830 44.680 5.990 46.090 ;
        RECT 6.180 45.275 6.440 45.945 ;
        RECT 6.195 44.885 6.425 45.275 ;
        RECT 6.620 44.680 6.780 46.090 ;
        RECT 6.985 45.505 7.215 45.885 ;
        RECT 6.970 44.835 7.230 45.505 ;
        RECT 7.410 44.680 7.570 46.090 ;
        RECT 7.760 45.275 8.020 45.945 ;
        RECT 7.775 44.885 8.005 45.275 ;
        RECT 8.200 44.680 8.360 46.090 ;
        RECT 8.565 45.505 8.795 45.885 ;
        RECT 8.550 44.835 8.810 45.505 ;
        RECT 8.990 44.680 9.150 46.090 ;
        RECT 9.340 45.275 9.600 45.945 ;
        RECT 9.355 44.885 9.585 45.275 ;
        RECT 9.780 44.680 9.940 46.090 ;
        RECT 10.145 45.505 10.375 45.885 ;
        RECT 10.130 44.835 10.390 45.505 ;
        RECT 10.570 44.680 10.730 46.090 ;
        RECT 10.920 45.275 11.180 45.945 ;
        RECT 10.935 44.885 11.165 45.275 ;
        RECT 11.360 44.680 11.520 46.090 ;
        RECT 11.725 45.505 11.955 45.885 ;
        RECT 11.710 44.835 11.970 45.505 ;
        RECT 12.150 44.680 12.310 46.090 ;
        RECT 12.500 45.275 12.760 45.945 ;
        RECT 12.515 44.885 12.745 45.275 ;
        RECT 12.940 44.680 13.100 46.090 ;
        RECT 13.305 45.505 13.535 45.885 ;
        RECT 13.290 44.835 13.550 45.505 ;
        RECT 13.730 44.680 13.890 46.090 ;
        RECT 14.080 45.275 14.340 45.945 ;
        RECT 14.095 44.885 14.325 45.275 ;
        RECT 14.520 44.680 14.680 46.090 ;
        RECT 14.885 45.505 15.115 45.885 ;
        RECT 14.870 44.835 15.130 45.505 ;
        RECT 15.310 44.680 15.470 46.090 ;
        RECT 15.660 45.275 15.920 45.945 ;
        RECT 15.675 44.885 15.905 45.275 ;
        RECT 16.100 44.680 16.260 46.090 ;
        RECT 16.465 45.505 16.695 45.885 ;
        RECT 16.450 44.835 16.710 45.505 ;
        RECT 16.890 44.680 17.050 46.090 ;
        RECT 17.240 45.275 17.500 45.945 ;
        RECT 17.255 44.885 17.485 45.275 ;
        RECT 17.680 44.680 17.840 46.090 ;
        RECT 18.045 45.505 18.275 45.885 ;
        RECT 18.030 44.835 18.290 45.505 ;
        RECT 18.470 44.680 18.630 46.090 ;
        RECT 18.820 45.275 19.080 45.945 ;
        RECT 18.835 44.885 19.065 45.275 ;
        RECT 2.525 44.660 3.775 44.680 ;
        RECT 4.105 44.660 4.565 44.680 ;
        RECT 4.895 44.660 5.355 44.680 ;
        RECT 5.685 44.660 6.145 44.680 ;
        RECT 6.475 44.660 6.935 44.680 ;
        RECT 7.265 44.660 7.725 44.680 ;
        RECT 8.055 44.660 8.515 44.680 ;
        RECT 8.845 44.660 9.305 44.680 ;
        RECT 9.635 44.660 10.095 44.680 ;
        RECT 10.425 44.660 10.885 44.680 ;
        RECT 11.215 44.660 11.675 44.680 ;
        RECT 12.005 44.660 12.465 44.680 ;
        RECT 12.795 44.660 13.255 44.680 ;
        RECT 13.585 44.660 14.045 44.680 ;
        RECT 14.375 44.660 14.835 44.680 ;
        RECT 15.165 44.660 15.625 44.680 ;
        RECT 15.955 44.660 16.415 44.680 ;
        RECT 16.745 44.660 17.205 44.680 ;
        RECT 17.535 44.660 17.995 44.680 ;
        RECT 18.325 44.660 18.785 44.680 ;
        RECT 2.525 44.475 18.785 44.660 ;
        RECT 2.525 44.450 3.775 44.475 ;
        RECT 4.105 44.450 4.565 44.475 ;
        RECT 4.895 44.450 5.355 44.475 ;
        RECT 5.685 44.450 6.145 44.475 ;
        RECT 6.475 44.450 6.935 44.475 ;
        RECT 7.265 44.450 7.725 44.475 ;
        RECT 8.055 44.450 8.515 44.475 ;
        RECT 8.845 44.450 9.305 44.475 ;
        RECT 9.635 44.450 10.095 44.475 ;
        RECT 10.425 44.450 10.885 44.475 ;
        RECT 11.215 44.450 11.675 44.475 ;
        RECT 12.005 44.450 12.465 44.475 ;
        RECT 12.795 44.450 13.255 44.475 ;
        RECT 13.585 44.450 14.045 44.475 ;
        RECT 14.375 44.450 14.835 44.475 ;
        RECT 15.165 44.450 15.625 44.475 ;
        RECT 15.955 44.450 16.415 44.475 ;
        RECT 16.745 44.450 17.205 44.475 ;
        RECT 17.535 44.450 17.995 44.475 ;
        RECT 18.325 44.450 18.785 44.475 ;
        RECT 2.525 44.140 2.760 44.450 ;
        RECT 3.460 44.140 3.620 44.450 ;
        RECT 4.250 44.140 4.410 44.450 ;
        RECT 5.040 44.140 5.200 44.450 ;
        RECT 5.830 44.140 5.990 44.450 ;
        RECT 6.620 44.140 6.780 44.450 ;
        RECT 7.410 44.140 7.570 44.450 ;
        RECT 8.200 44.140 8.360 44.450 ;
        RECT 8.990 44.140 9.150 44.450 ;
        RECT 9.780 44.140 9.940 44.450 ;
        RECT 10.570 44.140 10.730 44.450 ;
        RECT 11.360 44.140 11.520 44.450 ;
        RECT 12.150 44.140 12.310 44.450 ;
        RECT 12.940 44.140 13.100 44.450 ;
        RECT 13.730 44.140 13.890 44.450 ;
        RECT 14.520 44.140 14.680 44.450 ;
        RECT 15.310 44.140 15.470 44.450 ;
        RECT 16.100 44.140 16.260 44.450 ;
        RECT 16.890 44.140 17.050 44.450 ;
        RECT 17.680 44.140 17.840 44.450 ;
        RECT 18.470 44.140 18.630 44.450 ;
        RECT 2.525 44.120 3.775 44.140 ;
        RECT 4.105 44.120 4.565 44.140 ;
        RECT 4.895 44.120 5.355 44.140 ;
        RECT 5.685 44.120 6.145 44.140 ;
        RECT 6.475 44.120 6.935 44.140 ;
        RECT 7.265 44.120 7.725 44.140 ;
        RECT 8.055 44.120 8.515 44.140 ;
        RECT 8.845 44.120 9.305 44.140 ;
        RECT 9.635 44.120 10.095 44.140 ;
        RECT 10.425 44.120 10.885 44.140 ;
        RECT 11.215 44.120 11.675 44.140 ;
        RECT 12.005 44.120 12.465 44.140 ;
        RECT 12.795 44.120 13.255 44.140 ;
        RECT 13.585 44.120 14.045 44.140 ;
        RECT 14.375 44.120 14.835 44.140 ;
        RECT 15.165 44.120 15.625 44.140 ;
        RECT 15.955 44.120 16.415 44.140 ;
        RECT 16.745 44.120 17.205 44.140 ;
        RECT 17.535 44.120 17.995 44.140 ;
        RECT 18.325 44.120 18.785 44.140 ;
        RECT 2.525 43.935 18.825 44.120 ;
        RECT 2.525 43.910 3.775 43.935 ;
        RECT 4.105 43.910 4.565 43.935 ;
        RECT 4.895 43.910 5.355 43.935 ;
        RECT 5.685 43.910 6.145 43.935 ;
        RECT 6.475 43.910 6.935 43.935 ;
        RECT 7.265 43.910 7.725 43.935 ;
        RECT 8.055 43.910 8.515 43.935 ;
        RECT 8.845 43.910 9.305 43.935 ;
        RECT 9.635 43.910 10.095 43.935 ;
        RECT 10.425 43.910 10.885 43.935 ;
        RECT 11.215 43.910 11.675 43.935 ;
        RECT 12.005 43.910 12.465 43.935 ;
        RECT 12.795 43.910 13.255 43.935 ;
        RECT 13.585 43.910 14.045 43.935 ;
        RECT 14.375 43.910 14.835 43.935 ;
        RECT 15.165 43.910 15.625 43.935 ;
        RECT 15.955 43.910 16.415 43.935 ;
        RECT 16.745 43.910 17.205 43.935 ;
        RECT 17.535 43.910 17.995 43.935 ;
        RECT 18.325 43.910 18.785 43.935 ;
        RECT 2.525 42.500 2.760 43.910 ;
        RECT 3.020 43.095 3.280 43.765 ;
        RECT 3.035 42.705 3.265 43.095 ;
        RECT 3.460 42.500 3.620 43.910 ;
        RECT 3.825 43.325 4.055 43.705 ;
        RECT 3.810 42.655 4.070 43.325 ;
        RECT 4.250 42.500 4.410 43.910 ;
        RECT 4.600 43.095 4.860 43.765 ;
        RECT 4.615 42.705 4.845 43.095 ;
        RECT 5.040 42.500 5.200 43.910 ;
        RECT 5.405 43.325 5.635 43.705 ;
        RECT 5.390 42.655 5.650 43.325 ;
        RECT 5.830 42.500 5.990 43.910 ;
        RECT 6.180 43.095 6.440 43.765 ;
        RECT 6.195 42.705 6.425 43.095 ;
        RECT 6.620 42.500 6.780 43.910 ;
        RECT 6.985 43.325 7.215 43.705 ;
        RECT 6.970 42.655 7.230 43.325 ;
        RECT 7.410 42.500 7.570 43.910 ;
        RECT 7.760 43.095 8.020 43.765 ;
        RECT 7.775 42.705 8.005 43.095 ;
        RECT 8.200 42.500 8.360 43.910 ;
        RECT 8.565 43.325 8.795 43.705 ;
        RECT 8.550 42.655 8.810 43.325 ;
        RECT 8.990 42.500 9.150 43.910 ;
        RECT 9.340 43.095 9.600 43.765 ;
        RECT 9.355 42.705 9.585 43.095 ;
        RECT 9.780 42.500 9.940 43.910 ;
        RECT 10.145 43.325 10.375 43.705 ;
        RECT 10.130 42.655 10.390 43.325 ;
        RECT 10.570 42.500 10.730 43.910 ;
        RECT 10.920 43.095 11.180 43.765 ;
        RECT 10.935 42.705 11.165 43.095 ;
        RECT 11.360 42.500 11.520 43.910 ;
        RECT 11.725 43.325 11.955 43.705 ;
        RECT 11.710 42.655 11.970 43.325 ;
        RECT 12.150 42.500 12.310 43.910 ;
        RECT 12.500 43.095 12.760 43.765 ;
        RECT 12.515 42.705 12.745 43.095 ;
        RECT 12.940 42.500 13.100 43.910 ;
        RECT 13.305 43.325 13.535 43.705 ;
        RECT 13.290 42.655 13.550 43.325 ;
        RECT 13.730 42.500 13.890 43.910 ;
        RECT 14.080 43.095 14.340 43.765 ;
        RECT 14.095 42.705 14.325 43.095 ;
        RECT 14.520 42.500 14.680 43.910 ;
        RECT 14.885 43.325 15.115 43.705 ;
        RECT 14.870 42.655 15.130 43.325 ;
        RECT 15.310 42.500 15.470 43.910 ;
        RECT 15.660 43.095 15.920 43.765 ;
        RECT 15.675 42.705 15.905 43.095 ;
        RECT 16.100 42.500 16.260 43.910 ;
        RECT 16.465 43.325 16.695 43.705 ;
        RECT 16.450 42.655 16.710 43.325 ;
        RECT 16.890 42.500 17.050 43.910 ;
        RECT 17.240 43.095 17.500 43.765 ;
        RECT 17.255 42.705 17.485 43.095 ;
        RECT 17.680 42.500 17.840 43.910 ;
        RECT 18.045 43.325 18.275 43.705 ;
        RECT 18.030 42.655 18.290 43.325 ;
        RECT 18.470 42.500 18.630 43.910 ;
        RECT 18.820 43.095 19.080 43.765 ;
        RECT 18.835 42.705 19.065 43.095 ;
        RECT 2.525 42.480 3.775 42.500 ;
        RECT 4.105 42.480 4.565 42.500 ;
        RECT 4.895 42.480 5.355 42.500 ;
        RECT 5.685 42.480 6.145 42.500 ;
        RECT 6.475 42.480 6.935 42.500 ;
        RECT 7.265 42.480 7.725 42.500 ;
        RECT 8.055 42.480 8.515 42.500 ;
        RECT 8.845 42.480 9.305 42.500 ;
        RECT 9.635 42.480 10.095 42.500 ;
        RECT 10.425 42.480 10.885 42.500 ;
        RECT 11.215 42.480 11.675 42.500 ;
        RECT 12.005 42.480 12.465 42.500 ;
        RECT 12.795 42.480 13.255 42.500 ;
        RECT 13.585 42.480 14.045 42.500 ;
        RECT 14.375 42.480 14.835 42.500 ;
        RECT 15.165 42.480 15.625 42.500 ;
        RECT 15.955 42.480 16.415 42.500 ;
        RECT 16.745 42.480 17.205 42.500 ;
        RECT 17.535 42.480 17.995 42.500 ;
        RECT 18.325 42.480 18.785 42.500 ;
        RECT 2.525 42.295 18.785 42.480 ;
        RECT 2.525 42.270 3.775 42.295 ;
        RECT 4.105 42.270 4.565 42.295 ;
        RECT 4.895 42.270 5.355 42.295 ;
        RECT 5.685 42.270 6.145 42.295 ;
        RECT 6.475 42.270 6.935 42.295 ;
        RECT 7.265 42.270 7.725 42.295 ;
        RECT 8.055 42.270 8.515 42.295 ;
        RECT 8.845 42.270 9.305 42.295 ;
        RECT 9.635 42.270 10.095 42.295 ;
        RECT 10.425 42.270 10.885 42.295 ;
        RECT 11.215 42.270 11.675 42.295 ;
        RECT 12.005 42.270 12.465 42.295 ;
        RECT 12.795 42.270 13.255 42.295 ;
        RECT 13.585 42.270 14.045 42.295 ;
        RECT 14.375 42.270 14.835 42.295 ;
        RECT 15.165 42.270 15.625 42.295 ;
        RECT 15.955 42.270 16.415 42.295 ;
        RECT 16.745 42.270 17.205 42.295 ;
        RECT 17.535 42.270 17.995 42.295 ;
        RECT 18.325 42.270 18.785 42.295 ;
        RECT 2.525 41.960 2.760 42.270 ;
        RECT 3.460 41.960 3.620 42.270 ;
        RECT 4.250 41.960 4.410 42.270 ;
        RECT 5.040 41.960 5.200 42.270 ;
        RECT 5.830 41.960 5.990 42.270 ;
        RECT 6.620 41.960 6.780 42.270 ;
        RECT 7.410 41.960 7.570 42.270 ;
        RECT 8.200 41.960 8.360 42.270 ;
        RECT 8.990 41.960 9.150 42.270 ;
        RECT 9.780 41.960 9.940 42.270 ;
        RECT 10.570 41.960 10.730 42.270 ;
        RECT 11.360 41.960 11.520 42.270 ;
        RECT 12.150 41.960 12.310 42.270 ;
        RECT 12.940 41.960 13.100 42.270 ;
        RECT 13.730 41.960 13.890 42.270 ;
        RECT 14.520 41.960 14.680 42.270 ;
        RECT 15.310 41.960 15.470 42.270 ;
        RECT 16.100 41.960 16.260 42.270 ;
        RECT 16.890 41.960 17.050 42.270 ;
        RECT 17.680 41.960 17.840 42.270 ;
        RECT 18.470 41.960 18.630 42.270 ;
        RECT 2.525 41.940 3.775 41.960 ;
        RECT 4.105 41.940 4.565 41.960 ;
        RECT 4.895 41.940 5.355 41.960 ;
        RECT 5.685 41.940 6.145 41.960 ;
        RECT 6.475 41.940 6.935 41.960 ;
        RECT 7.265 41.940 7.725 41.960 ;
        RECT 8.055 41.940 8.515 41.960 ;
        RECT 8.845 41.940 9.305 41.960 ;
        RECT 9.635 41.940 10.095 41.960 ;
        RECT 10.425 41.940 10.885 41.960 ;
        RECT 11.215 41.940 11.675 41.960 ;
        RECT 12.005 41.940 12.465 41.960 ;
        RECT 12.795 41.940 13.255 41.960 ;
        RECT 13.585 41.940 14.045 41.960 ;
        RECT 14.375 41.940 14.835 41.960 ;
        RECT 15.165 41.940 15.625 41.960 ;
        RECT 15.955 41.940 16.415 41.960 ;
        RECT 16.745 41.940 17.205 41.960 ;
        RECT 17.535 41.940 17.995 41.960 ;
        RECT 18.325 41.940 18.785 41.960 ;
        RECT 2.525 41.755 18.825 41.940 ;
        RECT 2.525 41.730 3.775 41.755 ;
        RECT 4.105 41.730 4.565 41.755 ;
        RECT 4.895 41.730 5.355 41.755 ;
        RECT 5.685 41.730 6.145 41.755 ;
        RECT 6.475 41.730 6.935 41.755 ;
        RECT 7.265 41.730 7.725 41.755 ;
        RECT 8.055 41.730 8.515 41.755 ;
        RECT 8.845 41.730 9.305 41.755 ;
        RECT 9.635 41.730 10.095 41.755 ;
        RECT 10.425 41.730 10.885 41.755 ;
        RECT 11.215 41.730 11.675 41.755 ;
        RECT 12.005 41.730 12.465 41.755 ;
        RECT 12.795 41.730 13.255 41.755 ;
        RECT 13.585 41.730 14.045 41.755 ;
        RECT 14.375 41.730 14.835 41.755 ;
        RECT 15.165 41.730 15.625 41.755 ;
        RECT 15.955 41.730 16.415 41.755 ;
        RECT 16.745 41.730 17.205 41.755 ;
        RECT 17.535 41.730 17.995 41.755 ;
        RECT 18.325 41.730 18.785 41.755 ;
        RECT 2.525 40.320 2.760 41.730 ;
        RECT 3.020 40.915 3.280 41.585 ;
        RECT 3.035 40.525 3.265 40.915 ;
        RECT 3.460 40.320 3.620 41.730 ;
        RECT 3.825 41.145 4.055 41.525 ;
        RECT 3.810 40.475 4.070 41.145 ;
        RECT 4.250 40.320 4.410 41.730 ;
        RECT 4.600 40.915 4.860 41.585 ;
        RECT 4.615 40.525 4.845 40.915 ;
        RECT 5.040 40.320 5.200 41.730 ;
        RECT 5.405 41.145 5.635 41.525 ;
        RECT 5.390 40.475 5.650 41.145 ;
        RECT 5.830 40.320 5.990 41.730 ;
        RECT 6.180 40.915 6.440 41.585 ;
        RECT 6.195 40.525 6.425 40.915 ;
        RECT 6.620 40.320 6.780 41.730 ;
        RECT 6.985 41.145 7.215 41.525 ;
        RECT 6.970 40.475 7.230 41.145 ;
        RECT 7.410 40.320 7.570 41.730 ;
        RECT 7.760 40.915 8.020 41.585 ;
        RECT 7.775 40.525 8.005 40.915 ;
        RECT 8.200 40.320 8.360 41.730 ;
        RECT 8.565 41.145 8.795 41.525 ;
        RECT 8.550 40.475 8.810 41.145 ;
        RECT 8.990 40.320 9.150 41.730 ;
        RECT 9.340 40.915 9.600 41.585 ;
        RECT 9.355 40.525 9.585 40.915 ;
        RECT 9.780 40.320 9.940 41.730 ;
        RECT 10.145 41.145 10.375 41.525 ;
        RECT 10.130 40.475 10.390 41.145 ;
        RECT 10.570 40.320 10.730 41.730 ;
        RECT 10.920 40.915 11.180 41.585 ;
        RECT 10.935 40.525 11.165 40.915 ;
        RECT 11.360 40.320 11.520 41.730 ;
        RECT 11.725 41.145 11.955 41.525 ;
        RECT 11.710 40.475 11.970 41.145 ;
        RECT 12.150 40.320 12.310 41.730 ;
        RECT 12.500 40.915 12.760 41.585 ;
        RECT 12.515 40.525 12.745 40.915 ;
        RECT 12.940 40.320 13.100 41.730 ;
        RECT 13.305 41.145 13.535 41.525 ;
        RECT 13.290 40.475 13.550 41.145 ;
        RECT 13.730 40.320 13.890 41.730 ;
        RECT 14.080 40.915 14.340 41.585 ;
        RECT 14.095 40.525 14.325 40.915 ;
        RECT 14.520 40.320 14.680 41.730 ;
        RECT 14.885 41.145 15.115 41.525 ;
        RECT 14.870 40.475 15.130 41.145 ;
        RECT 15.310 40.320 15.470 41.730 ;
        RECT 15.660 40.915 15.920 41.585 ;
        RECT 15.675 40.525 15.905 40.915 ;
        RECT 16.100 40.320 16.260 41.730 ;
        RECT 16.465 41.145 16.695 41.525 ;
        RECT 16.450 40.475 16.710 41.145 ;
        RECT 16.890 40.320 17.050 41.730 ;
        RECT 17.240 40.915 17.500 41.585 ;
        RECT 17.255 40.525 17.485 40.915 ;
        RECT 17.680 40.320 17.840 41.730 ;
        RECT 18.045 41.145 18.275 41.525 ;
        RECT 18.030 40.475 18.290 41.145 ;
        RECT 18.470 40.320 18.630 41.730 ;
        RECT 18.820 40.915 19.080 41.585 ;
        RECT 18.835 40.525 19.065 40.915 ;
        RECT 2.525 40.300 3.775 40.320 ;
        RECT 4.105 40.300 4.565 40.320 ;
        RECT 4.895 40.300 5.355 40.320 ;
        RECT 5.685 40.300 6.145 40.320 ;
        RECT 6.475 40.300 6.935 40.320 ;
        RECT 7.265 40.300 7.725 40.320 ;
        RECT 8.055 40.300 8.515 40.320 ;
        RECT 8.845 40.300 9.305 40.320 ;
        RECT 9.635 40.300 10.095 40.320 ;
        RECT 10.425 40.300 10.885 40.320 ;
        RECT 11.215 40.300 11.675 40.320 ;
        RECT 12.005 40.300 12.465 40.320 ;
        RECT 12.795 40.300 13.255 40.320 ;
        RECT 13.585 40.300 14.045 40.320 ;
        RECT 14.375 40.300 14.835 40.320 ;
        RECT 15.165 40.300 15.625 40.320 ;
        RECT 15.955 40.300 16.415 40.320 ;
        RECT 16.745 40.300 17.205 40.320 ;
        RECT 17.535 40.300 17.995 40.320 ;
        RECT 18.325 40.300 18.785 40.320 ;
        RECT 2.525 40.115 18.785 40.300 ;
        RECT 2.525 40.090 3.775 40.115 ;
        RECT 4.105 40.090 4.565 40.115 ;
        RECT 4.895 40.090 5.355 40.115 ;
        RECT 5.685 40.090 6.145 40.115 ;
        RECT 6.475 40.090 6.935 40.115 ;
        RECT 7.265 40.090 7.725 40.115 ;
        RECT 8.055 40.090 8.515 40.115 ;
        RECT 8.845 40.090 9.305 40.115 ;
        RECT 9.635 40.090 10.095 40.115 ;
        RECT 10.425 40.090 10.885 40.115 ;
        RECT 11.215 40.090 11.675 40.115 ;
        RECT 12.005 40.090 12.465 40.115 ;
        RECT 12.795 40.090 13.255 40.115 ;
        RECT 13.585 40.090 14.045 40.115 ;
        RECT 14.375 40.090 14.835 40.115 ;
        RECT 15.165 40.090 15.625 40.115 ;
        RECT 15.955 40.090 16.415 40.115 ;
        RECT 16.745 40.090 17.205 40.115 ;
        RECT 17.535 40.090 17.995 40.115 ;
        RECT 18.325 40.090 18.785 40.115 ;
        RECT 2.525 39.780 2.760 40.090 ;
        RECT 3.460 39.780 3.620 40.090 ;
        RECT 4.250 39.780 4.410 40.090 ;
        RECT 5.040 39.780 5.200 40.090 ;
        RECT 5.830 39.780 5.990 40.090 ;
        RECT 6.620 39.780 6.780 40.090 ;
        RECT 7.410 39.780 7.570 40.090 ;
        RECT 8.200 39.780 8.360 40.090 ;
        RECT 8.990 39.780 9.150 40.090 ;
        RECT 9.780 39.780 9.940 40.090 ;
        RECT 10.570 39.780 10.730 40.090 ;
        RECT 11.360 39.780 11.520 40.090 ;
        RECT 12.150 39.780 12.310 40.090 ;
        RECT 12.940 39.780 13.100 40.090 ;
        RECT 13.730 39.780 13.890 40.090 ;
        RECT 14.520 39.780 14.680 40.090 ;
        RECT 15.310 39.780 15.470 40.090 ;
        RECT 16.100 39.780 16.260 40.090 ;
        RECT 16.890 39.780 17.050 40.090 ;
        RECT 17.680 39.780 17.840 40.090 ;
        RECT 18.470 39.780 18.630 40.090 ;
        RECT 2.525 39.760 3.775 39.780 ;
        RECT 4.105 39.760 4.565 39.780 ;
        RECT 4.895 39.760 5.355 39.780 ;
        RECT 5.685 39.760 6.145 39.780 ;
        RECT 6.475 39.760 6.935 39.780 ;
        RECT 7.265 39.760 7.725 39.780 ;
        RECT 8.055 39.760 8.515 39.780 ;
        RECT 8.845 39.760 9.305 39.780 ;
        RECT 9.635 39.760 10.095 39.780 ;
        RECT 10.425 39.760 10.885 39.780 ;
        RECT 11.215 39.760 11.675 39.780 ;
        RECT 12.005 39.760 12.465 39.780 ;
        RECT 12.795 39.760 13.255 39.780 ;
        RECT 13.585 39.760 14.045 39.780 ;
        RECT 14.375 39.760 14.835 39.780 ;
        RECT 15.165 39.760 15.625 39.780 ;
        RECT 15.955 39.760 16.415 39.780 ;
        RECT 16.745 39.760 17.205 39.780 ;
        RECT 17.535 39.760 17.995 39.780 ;
        RECT 18.325 39.760 18.785 39.780 ;
        RECT 2.525 39.575 18.825 39.760 ;
        RECT 2.525 39.550 3.775 39.575 ;
        RECT 4.105 39.550 4.565 39.575 ;
        RECT 4.895 39.550 5.355 39.575 ;
        RECT 5.685 39.550 6.145 39.575 ;
        RECT 6.475 39.550 6.935 39.575 ;
        RECT 7.265 39.550 7.725 39.575 ;
        RECT 8.055 39.550 8.515 39.575 ;
        RECT 8.845 39.550 9.305 39.575 ;
        RECT 9.635 39.550 10.095 39.575 ;
        RECT 10.425 39.550 10.885 39.575 ;
        RECT 11.215 39.550 11.675 39.575 ;
        RECT 12.005 39.550 12.465 39.575 ;
        RECT 12.795 39.550 13.255 39.575 ;
        RECT 13.585 39.550 14.045 39.575 ;
        RECT 14.375 39.550 14.835 39.575 ;
        RECT 15.165 39.550 15.625 39.575 ;
        RECT 15.955 39.550 16.415 39.575 ;
        RECT 16.745 39.550 17.205 39.575 ;
        RECT 17.535 39.550 17.995 39.575 ;
        RECT 18.325 39.550 18.785 39.575 ;
        RECT 2.525 38.140 2.760 39.550 ;
        RECT 3.020 38.735 3.280 39.405 ;
        RECT 3.035 38.345 3.265 38.735 ;
        RECT 3.460 38.140 3.620 39.550 ;
        RECT 3.825 38.965 4.055 39.345 ;
        RECT 3.810 38.295 4.070 38.965 ;
        RECT 4.250 38.140 4.410 39.550 ;
        RECT 4.600 38.735 4.860 39.405 ;
        RECT 4.615 38.345 4.845 38.735 ;
        RECT 5.040 38.140 5.200 39.550 ;
        RECT 5.405 38.965 5.635 39.345 ;
        RECT 5.390 38.295 5.650 38.965 ;
        RECT 5.830 38.140 5.990 39.550 ;
        RECT 6.180 38.735 6.440 39.405 ;
        RECT 6.195 38.345 6.425 38.735 ;
        RECT 6.620 38.140 6.780 39.550 ;
        RECT 6.985 38.965 7.215 39.345 ;
        RECT 6.970 38.295 7.230 38.965 ;
        RECT 7.410 38.140 7.570 39.550 ;
        RECT 7.760 38.735 8.020 39.405 ;
        RECT 7.775 38.345 8.005 38.735 ;
        RECT 8.200 38.140 8.360 39.550 ;
        RECT 8.565 38.965 8.795 39.345 ;
        RECT 8.550 38.295 8.810 38.965 ;
        RECT 8.990 38.140 9.150 39.550 ;
        RECT 9.340 38.735 9.600 39.405 ;
        RECT 9.355 38.345 9.585 38.735 ;
        RECT 9.780 38.140 9.940 39.550 ;
        RECT 10.145 38.965 10.375 39.345 ;
        RECT 10.130 38.295 10.390 38.965 ;
        RECT 10.570 38.140 10.730 39.550 ;
        RECT 10.920 38.735 11.180 39.405 ;
        RECT 10.935 38.345 11.165 38.735 ;
        RECT 11.360 38.140 11.520 39.550 ;
        RECT 11.725 38.965 11.955 39.345 ;
        RECT 11.710 38.295 11.970 38.965 ;
        RECT 12.150 38.140 12.310 39.550 ;
        RECT 12.500 38.735 12.760 39.405 ;
        RECT 12.515 38.345 12.745 38.735 ;
        RECT 12.940 38.140 13.100 39.550 ;
        RECT 13.305 38.965 13.535 39.345 ;
        RECT 13.290 38.295 13.550 38.965 ;
        RECT 13.730 38.140 13.890 39.550 ;
        RECT 14.080 38.735 14.340 39.405 ;
        RECT 14.095 38.345 14.325 38.735 ;
        RECT 14.520 38.140 14.680 39.550 ;
        RECT 14.885 38.965 15.115 39.345 ;
        RECT 14.870 38.295 15.130 38.965 ;
        RECT 15.310 38.140 15.470 39.550 ;
        RECT 15.660 38.735 15.920 39.405 ;
        RECT 15.675 38.345 15.905 38.735 ;
        RECT 16.100 38.140 16.260 39.550 ;
        RECT 16.465 38.965 16.695 39.345 ;
        RECT 16.450 38.295 16.710 38.965 ;
        RECT 16.890 38.140 17.050 39.550 ;
        RECT 17.240 38.735 17.500 39.405 ;
        RECT 17.255 38.345 17.485 38.735 ;
        RECT 17.680 38.140 17.840 39.550 ;
        RECT 18.045 38.965 18.275 39.345 ;
        RECT 18.030 38.295 18.290 38.965 ;
        RECT 18.470 38.140 18.630 39.550 ;
        RECT 18.820 38.735 19.080 39.405 ;
        RECT 18.835 38.345 19.065 38.735 ;
        RECT 2.525 38.120 3.775 38.140 ;
        RECT 4.105 38.120 4.565 38.140 ;
        RECT 4.895 38.120 5.355 38.140 ;
        RECT 5.685 38.120 6.145 38.140 ;
        RECT 6.475 38.120 6.935 38.140 ;
        RECT 7.265 38.120 7.725 38.140 ;
        RECT 8.055 38.120 8.515 38.140 ;
        RECT 8.845 38.120 9.305 38.140 ;
        RECT 9.635 38.120 10.095 38.140 ;
        RECT 10.425 38.120 10.885 38.140 ;
        RECT 11.215 38.120 11.675 38.140 ;
        RECT 12.005 38.120 12.465 38.140 ;
        RECT 12.795 38.120 13.255 38.140 ;
        RECT 13.585 38.120 14.045 38.140 ;
        RECT 14.375 38.120 14.835 38.140 ;
        RECT 15.165 38.120 15.625 38.140 ;
        RECT 15.955 38.120 16.415 38.140 ;
        RECT 16.745 38.120 17.205 38.140 ;
        RECT 17.535 38.120 17.995 38.140 ;
        RECT 18.325 38.120 18.785 38.140 ;
        RECT 2.525 37.935 18.785 38.120 ;
        RECT 2.525 37.910 3.775 37.935 ;
        RECT 4.105 37.910 4.565 37.935 ;
        RECT 4.895 37.910 5.355 37.935 ;
        RECT 5.685 37.910 6.145 37.935 ;
        RECT 6.475 37.910 6.935 37.935 ;
        RECT 7.265 37.910 7.725 37.935 ;
        RECT 8.055 37.910 8.515 37.935 ;
        RECT 8.845 37.910 9.305 37.935 ;
        RECT 9.635 37.910 10.095 37.935 ;
        RECT 10.425 37.910 10.885 37.935 ;
        RECT 11.215 37.910 11.675 37.935 ;
        RECT 12.005 37.910 12.465 37.935 ;
        RECT 12.795 37.910 13.255 37.935 ;
        RECT 13.585 37.910 14.045 37.935 ;
        RECT 14.375 37.910 14.835 37.935 ;
        RECT 15.165 37.910 15.625 37.935 ;
        RECT 15.955 37.910 16.415 37.935 ;
        RECT 16.745 37.910 17.205 37.935 ;
        RECT 17.535 37.910 17.995 37.935 ;
        RECT 18.325 37.910 18.785 37.935 ;
        RECT 2.525 37.600 2.760 37.910 ;
        RECT 3.460 37.600 3.620 37.910 ;
        RECT 4.250 37.600 4.410 37.910 ;
        RECT 5.040 37.600 5.200 37.910 ;
        RECT 5.830 37.600 5.990 37.910 ;
        RECT 6.620 37.600 6.780 37.910 ;
        RECT 7.410 37.600 7.570 37.910 ;
        RECT 8.200 37.600 8.360 37.910 ;
        RECT 8.990 37.600 9.150 37.910 ;
        RECT 9.780 37.600 9.940 37.910 ;
        RECT 10.570 37.600 10.730 37.910 ;
        RECT 11.360 37.600 11.520 37.910 ;
        RECT 12.150 37.600 12.310 37.910 ;
        RECT 12.940 37.600 13.100 37.910 ;
        RECT 13.730 37.600 13.890 37.910 ;
        RECT 14.520 37.600 14.680 37.910 ;
        RECT 15.310 37.600 15.470 37.910 ;
        RECT 16.100 37.600 16.260 37.910 ;
        RECT 16.890 37.600 17.050 37.910 ;
        RECT 17.680 37.600 17.840 37.910 ;
        RECT 18.470 37.600 18.630 37.910 ;
        RECT 2.525 37.580 3.775 37.600 ;
        RECT 4.105 37.580 4.565 37.600 ;
        RECT 4.895 37.580 5.355 37.600 ;
        RECT 5.685 37.580 6.145 37.600 ;
        RECT 6.475 37.580 6.935 37.600 ;
        RECT 7.265 37.580 7.725 37.600 ;
        RECT 8.055 37.580 8.515 37.600 ;
        RECT 8.845 37.580 9.305 37.600 ;
        RECT 9.635 37.580 10.095 37.600 ;
        RECT 10.425 37.580 10.885 37.600 ;
        RECT 11.215 37.580 11.675 37.600 ;
        RECT 12.005 37.580 12.465 37.600 ;
        RECT 12.795 37.580 13.255 37.600 ;
        RECT 13.585 37.580 14.045 37.600 ;
        RECT 14.375 37.580 14.835 37.600 ;
        RECT 15.165 37.580 15.625 37.600 ;
        RECT 15.955 37.580 16.415 37.600 ;
        RECT 16.745 37.580 17.205 37.600 ;
        RECT 17.535 37.580 17.995 37.600 ;
        RECT 18.325 37.580 18.785 37.600 ;
        RECT 2.525 37.395 18.825 37.580 ;
        RECT 2.525 37.370 3.775 37.395 ;
        RECT 4.105 37.370 4.565 37.395 ;
        RECT 4.895 37.370 5.355 37.395 ;
        RECT 5.685 37.370 6.145 37.395 ;
        RECT 6.475 37.370 6.935 37.395 ;
        RECT 7.265 37.370 7.725 37.395 ;
        RECT 8.055 37.370 8.515 37.395 ;
        RECT 8.845 37.370 9.305 37.395 ;
        RECT 9.635 37.370 10.095 37.395 ;
        RECT 10.425 37.370 10.885 37.395 ;
        RECT 11.215 37.370 11.675 37.395 ;
        RECT 12.005 37.370 12.465 37.395 ;
        RECT 12.795 37.370 13.255 37.395 ;
        RECT 13.585 37.370 14.045 37.395 ;
        RECT 14.375 37.370 14.835 37.395 ;
        RECT 15.165 37.370 15.625 37.395 ;
        RECT 15.955 37.370 16.415 37.395 ;
        RECT 16.745 37.370 17.205 37.395 ;
        RECT 17.535 37.370 17.995 37.395 ;
        RECT 18.325 37.370 18.785 37.395 ;
        RECT 2.525 35.960 2.760 37.370 ;
        RECT 3.020 36.555 3.280 37.225 ;
        RECT 3.035 36.165 3.265 36.555 ;
        RECT 3.460 35.960 3.620 37.370 ;
        RECT 3.825 36.785 4.055 37.165 ;
        RECT 3.810 36.115 4.070 36.785 ;
        RECT 4.250 35.960 4.410 37.370 ;
        RECT 4.600 36.555 4.860 37.225 ;
        RECT 4.615 36.165 4.845 36.555 ;
        RECT 5.040 35.960 5.200 37.370 ;
        RECT 5.405 36.785 5.635 37.165 ;
        RECT 5.390 36.115 5.650 36.785 ;
        RECT 5.830 35.960 5.990 37.370 ;
        RECT 6.180 36.555 6.440 37.225 ;
        RECT 6.195 36.165 6.425 36.555 ;
        RECT 6.620 35.960 6.780 37.370 ;
        RECT 6.985 36.785 7.215 37.165 ;
        RECT 6.970 36.115 7.230 36.785 ;
        RECT 7.410 35.960 7.570 37.370 ;
        RECT 7.760 36.555 8.020 37.225 ;
        RECT 7.775 36.165 8.005 36.555 ;
        RECT 8.200 35.960 8.360 37.370 ;
        RECT 8.565 36.785 8.795 37.165 ;
        RECT 8.550 36.115 8.810 36.785 ;
        RECT 8.990 35.960 9.150 37.370 ;
        RECT 9.340 36.555 9.600 37.225 ;
        RECT 9.355 36.165 9.585 36.555 ;
        RECT 9.780 35.960 9.940 37.370 ;
        RECT 10.145 36.785 10.375 37.165 ;
        RECT 10.130 36.115 10.390 36.785 ;
        RECT 10.570 35.960 10.730 37.370 ;
        RECT 10.920 36.555 11.180 37.225 ;
        RECT 10.935 36.165 11.165 36.555 ;
        RECT 11.360 35.960 11.520 37.370 ;
        RECT 11.725 36.785 11.955 37.165 ;
        RECT 11.710 36.115 11.970 36.785 ;
        RECT 12.150 35.960 12.310 37.370 ;
        RECT 12.500 36.555 12.760 37.225 ;
        RECT 12.515 36.165 12.745 36.555 ;
        RECT 12.940 35.960 13.100 37.370 ;
        RECT 13.305 36.785 13.535 37.165 ;
        RECT 13.290 36.115 13.550 36.785 ;
        RECT 13.730 35.960 13.890 37.370 ;
        RECT 14.080 36.555 14.340 37.225 ;
        RECT 14.095 36.165 14.325 36.555 ;
        RECT 14.520 35.960 14.680 37.370 ;
        RECT 14.885 36.785 15.115 37.165 ;
        RECT 14.870 36.115 15.130 36.785 ;
        RECT 15.310 35.960 15.470 37.370 ;
        RECT 15.660 36.555 15.920 37.225 ;
        RECT 15.675 36.165 15.905 36.555 ;
        RECT 16.100 35.960 16.260 37.370 ;
        RECT 16.465 36.785 16.695 37.165 ;
        RECT 16.450 36.115 16.710 36.785 ;
        RECT 16.890 35.960 17.050 37.370 ;
        RECT 17.240 36.555 17.500 37.225 ;
        RECT 17.255 36.165 17.485 36.555 ;
        RECT 17.680 35.960 17.840 37.370 ;
        RECT 18.045 36.785 18.275 37.165 ;
        RECT 18.030 36.115 18.290 36.785 ;
        RECT 18.470 35.960 18.630 37.370 ;
        RECT 18.820 36.555 19.080 37.225 ;
        RECT 18.835 36.165 19.065 36.555 ;
        RECT 2.525 35.940 3.775 35.960 ;
        RECT 4.105 35.940 4.565 35.960 ;
        RECT 4.895 35.940 5.355 35.960 ;
        RECT 5.685 35.940 6.145 35.960 ;
        RECT 6.475 35.940 6.935 35.960 ;
        RECT 7.265 35.940 7.725 35.960 ;
        RECT 8.055 35.940 8.515 35.960 ;
        RECT 8.845 35.940 9.305 35.960 ;
        RECT 9.635 35.940 10.095 35.960 ;
        RECT 10.425 35.940 10.885 35.960 ;
        RECT 11.215 35.940 11.675 35.960 ;
        RECT 12.005 35.940 12.465 35.960 ;
        RECT 12.795 35.940 13.255 35.960 ;
        RECT 13.585 35.940 14.045 35.960 ;
        RECT 14.375 35.940 14.835 35.960 ;
        RECT 15.165 35.940 15.625 35.960 ;
        RECT 15.955 35.940 16.415 35.960 ;
        RECT 16.745 35.940 17.205 35.960 ;
        RECT 17.535 35.940 17.995 35.960 ;
        RECT 18.325 35.940 18.785 35.960 ;
        RECT 2.525 35.755 18.785 35.940 ;
        RECT 2.525 35.730 3.775 35.755 ;
        RECT 4.105 35.730 4.565 35.755 ;
        RECT 4.895 35.730 5.355 35.755 ;
        RECT 5.685 35.730 6.145 35.755 ;
        RECT 6.475 35.730 6.935 35.755 ;
        RECT 7.265 35.730 7.725 35.755 ;
        RECT 8.055 35.730 8.515 35.755 ;
        RECT 8.845 35.730 9.305 35.755 ;
        RECT 9.635 35.730 10.095 35.755 ;
        RECT 10.425 35.730 10.885 35.755 ;
        RECT 11.215 35.730 11.675 35.755 ;
        RECT 12.005 35.730 12.465 35.755 ;
        RECT 12.795 35.730 13.255 35.755 ;
        RECT 13.585 35.730 14.045 35.755 ;
        RECT 14.375 35.730 14.835 35.755 ;
        RECT 15.165 35.730 15.625 35.755 ;
        RECT 15.955 35.730 16.415 35.755 ;
        RECT 16.745 35.730 17.205 35.755 ;
        RECT 17.535 35.730 17.995 35.755 ;
        RECT 18.325 35.730 18.785 35.755 ;
        RECT 2.525 35.420 2.760 35.730 ;
        RECT 3.460 35.420 3.620 35.730 ;
        RECT 4.250 35.420 4.410 35.730 ;
        RECT 5.040 35.420 5.200 35.730 ;
        RECT 5.830 35.420 5.990 35.730 ;
        RECT 6.620 35.420 6.780 35.730 ;
        RECT 7.410 35.420 7.570 35.730 ;
        RECT 8.200 35.420 8.360 35.730 ;
        RECT 8.990 35.420 9.150 35.730 ;
        RECT 9.780 35.420 9.940 35.730 ;
        RECT 10.570 35.420 10.730 35.730 ;
        RECT 11.360 35.420 11.520 35.730 ;
        RECT 12.150 35.420 12.310 35.730 ;
        RECT 12.940 35.420 13.100 35.730 ;
        RECT 13.730 35.420 13.890 35.730 ;
        RECT 14.520 35.420 14.680 35.730 ;
        RECT 15.310 35.420 15.470 35.730 ;
        RECT 16.100 35.420 16.260 35.730 ;
        RECT 16.890 35.420 17.050 35.730 ;
        RECT 17.680 35.420 17.840 35.730 ;
        RECT 18.470 35.420 18.630 35.730 ;
        RECT 2.525 35.400 3.775 35.420 ;
        RECT 4.105 35.400 4.565 35.420 ;
        RECT 4.895 35.400 5.355 35.420 ;
        RECT 5.685 35.400 6.145 35.420 ;
        RECT 6.475 35.400 6.935 35.420 ;
        RECT 7.265 35.400 7.725 35.420 ;
        RECT 8.055 35.400 8.515 35.420 ;
        RECT 8.845 35.400 9.305 35.420 ;
        RECT 9.635 35.400 10.095 35.420 ;
        RECT 10.425 35.400 10.885 35.420 ;
        RECT 11.215 35.400 11.675 35.420 ;
        RECT 12.005 35.400 12.465 35.420 ;
        RECT 12.795 35.400 13.255 35.420 ;
        RECT 13.585 35.400 14.045 35.420 ;
        RECT 14.375 35.400 14.835 35.420 ;
        RECT 15.165 35.400 15.625 35.420 ;
        RECT 15.955 35.400 16.415 35.420 ;
        RECT 16.745 35.400 17.205 35.420 ;
        RECT 17.535 35.400 17.995 35.420 ;
        RECT 18.325 35.400 18.785 35.420 ;
        RECT 2.525 35.215 18.825 35.400 ;
        RECT 2.525 35.190 3.775 35.215 ;
        RECT 4.105 35.190 4.565 35.215 ;
        RECT 4.895 35.190 5.355 35.215 ;
        RECT 5.685 35.190 6.145 35.215 ;
        RECT 6.475 35.190 6.935 35.215 ;
        RECT 7.265 35.190 7.725 35.215 ;
        RECT 8.055 35.190 8.515 35.215 ;
        RECT 8.845 35.190 9.305 35.215 ;
        RECT 9.635 35.190 10.095 35.215 ;
        RECT 10.425 35.190 10.885 35.215 ;
        RECT 11.215 35.190 11.675 35.215 ;
        RECT 12.005 35.190 12.465 35.215 ;
        RECT 12.795 35.190 13.255 35.215 ;
        RECT 13.585 35.190 14.045 35.215 ;
        RECT 14.375 35.190 14.835 35.215 ;
        RECT 15.165 35.190 15.625 35.215 ;
        RECT 15.955 35.190 16.415 35.215 ;
        RECT 16.745 35.190 17.205 35.215 ;
        RECT 17.535 35.190 17.995 35.215 ;
        RECT 18.325 35.190 18.785 35.215 ;
        RECT 2.525 33.780 2.760 35.190 ;
        RECT 3.020 34.375 3.280 35.045 ;
        RECT 3.035 33.985 3.265 34.375 ;
        RECT 3.460 33.780 3.620 35.190 ;
        RECT 3.825 34.605 4.055 34.985 ;
        RECT 3.810 33.935 4.070 34.605 ;
        RECT 4.250 33.780 4.410 35.190 ;
        RECT 4.600 34.375 4.860 35.045 ;
        RECT 4.615 33.985 4.845 34.375 ;
        RECT 5.040 33.780 5.200 35.190 ;
        RECT 5.405 34.605 5.635 34.985 ;
        RECT 5.390 33.935 5.650 34.605 ;
        RECT 5.830 33.780 5.990 35.190 ;
        RECT 6.180 34.375 6.440 35.045 ;
        RECT 6.195 33.985 6.425 34.375 ;
        RECT 6.620 33.780 6.780 35.190 ;
        RECT 6.985 34.605 7.215 34.985 ;
        RECT 6.970 33.935 7.230 34.605 ;
        RECT 7.410 33.780 7.570 35.190 ;
        RECT 7.760 34.375 8.020 35.045 ;
        RECT 7.775 33.985 8.005 34.375 ;
        RECT 8.200 33.780 8.360 35.190 ;
        RECT 8.565 34.605 8.795 34.985 ;
        RECT 8.550 33.935 8.810 34.605 ;
        RECT 8.990 33.780 9.150 35.190 ;
        RECT 9.340 34.375 9.600 35.045 ;
        RECT 9.355 33.985 9.585 34.375 ;
        RECT 9.780 33.780 9.940 35.190 ;
        RECT 10.145 34.605 10.375 34.985 ;
        RECT 10.130 33.935 10.390 34.605 ;
        RECT 10.570 33.780 10.730 35.190 ;
        RECT 10.920 34.375 11.180 35.045 ;
        RECT 10.935 33.985 11.165 34.375 ;
        RECT 11.360 33.780 11.520 35.190 ;
        RECT 11.725 34.605 11.955 34.985 ;
        RECT 11.710 33.935 11.970 34.605 ;
        RECT 12.150 33.780 12.310 35.190 ;
        RECT 12.500 34.375 12.760 35.045 ;
        RECT 12.515 33.985 12.745 34.375 ;
        RECT 12.940 33.780 13.100 35.190 ;
        RECT 13.305 34.605 13.535 34.985 ;
        RECT 13.290 33.935 13.550 34.605 ;
        RECT 13.730 33.780 13.890 35.190 ;
        RECT 14.080 34.375 14.340 35.045 ;
        RECT 14.095 33.985 14.325 34.375 ;
        RECT 14.520 33.780 14.680 35.190 ;
        RECT 14.885 34.605 15.115 34.985 ;
        RECT 14.870 33.935 15.130 34.605 ;
        RECT 15.310 33.780 15.470 35.190 ;
        RECT 15.660 34.375 15.920 35.045 ;
        RECT 15.675 33.985 15.905 34.375 ;
        RECT 16.100 33.780 16.260 35.190 ;
        RECT 16.465 34.605 16.695 34.985 ;
        RECT 16.450 33.935 16.710 34.605 ;
        RECT 16.890 33.780 17.050 35.190 ;
        RECT 17.240 34.375 17.500 35.045 ;
        RECT 17.255 33.985 17.485 34.375 ;
        RECT 17.680 33.780 17.840 35.190 ;
        RECT 18.045 34.605 18.275 34.985 ;
        RECT 18.030 33.935 18.290 34.605 ;
        RECT 18.470 33.780 18.630 35.190 ;
        RECT 18.820 34.375 19.080 35.045 ;
        RECT 18.835 33.985 19.065 34.375 ;
        RECT 2.525 33.760 3.775 33.780 ;
        RECT 4.105 33.760 4.565 33.780 ;
        RECT 4.895 33.760 5.355 33.780 ;
        RECT 5.685 33.760 6.145 33.780 ;
        RECT 6.475 33.760 6.935 33.780 ;
        RECT 7.265 33.760 7.725 33.780 ;
        RECT 8.055 33.760 8.515 33.780 ;
        RECT 8.845 33.760 9.305 33.780 ;
        RECT 9.635 33.760 10.095 33.780 ;
        RECT 10.425 33.760 10.885 33.780 ;
        RECT 11.215 33.760 11.675 33.780 ;
        RECT 12.005 33.760 12.465 33.780 ;
        RECT 12.795 33.760 13.255 33.780 ;
        RECT 13.585 33.760 14.045 33.780 ;
        RECT 14.375 33.760 14.835 33.780 ;
        RECT 15.165 33.760 15.625 33.780 ;
        RECT 15.955 33.760 16.415 33.780 ;
        RECT 16.745 33.760 17.205 33.780 ;
        RECT 17.535 33.760 17.995 33.780 ;
        RECT 18.325 33.760 18.785 33.780 ;
        RECT 2.525 33.575 18.785 33.760 ;
        RECT 2.525 33.550 3.775 33.575 ;
        RECT 4.105 33.550 4.565 33.575 ;
        RECT 4.895 33.550 5.355 33.575 ;
        RECT 5.685 33.550 6.145 33.575 ;
        RECT 6.475 33.550 6.935 33.575 ;
        RECT 7.265 33.550 7.725 33.575 ;
        RECT 8.055 33.550 8.515 33.575 ;
        RECT 8.845 33.550 9.305 33.575 ;
        RECT 9.635 33.550 10.095 33.575 ;
        RECT 10.425 33.550 10.885 33.575 ;
        RECT 11.215 33.550 11.675 33.575 ;
        RECT 12.005 33.550 12.465 33.575 ;
        RECT 12.795 33.550 13.255 33.575 ;
        RECT 13.585 33.550 14.045 33.575 ;
        RECT 14.375 33.550 14.835 33.575 ;
        RECT 15.165 33.550 15.625 33.575 ;
        RECT 15.955 33.550 16.415 33.575 ;
        RECT 16.745 33.550 17.205 33.575 ;
        RECT 17.535 33.550 17.995 33.575 ;
        RECT 18.325 33.550 18.785 33.575 ;
        RECT 2.525 33.240 2.760 33.550 ;
        RECT 3.460 33.240 3.620 33.550 ;
        RECT 4.250 33.240 4.410 33.550 ;
        RECT 5.040 33.240 5.200 33.550 ;
        RECT 5.830 33.240 5.990 33.550 ;
        RECT 6.620 33.240 6.780 33.550 ;
        RECT 7.410 33.240 7.570 33.550 ;
        RECT 8.200 33.240 8.360 33.550 ;
        RECT 8.990 33.240 9.150 33.550 ;
        RECT 9.780 33.240 9.940 33.550 ;
        RECT 10.570 33.240 10.730 33.550 ;
        RECT 11.360 33.240 11.520 33.550 ;
        RECT 12.150 33.240 12.310 33.550 ;
        RECT 12.940 33.240 13.100 33.550 ;
        RECT 13.730 33.240 13.890 33.550 ;
        RECT 14.520 33.240 14.680 33.550 ;
        RECT 15.310 33.240 15.470 33.550 ;
        RECT 16.100 33.240 16.260 33.550 ;
        RECT 16.890 33.240 17.050 33.550 ;
        RECT 17.680 33.240 17.840 33.550 ;
        RECT 18.470 33.240 18.630 33.550 ;
        RECT 2.525 33.220 3.775 33.240 ;
        RECT 4.105 33.220 4.565 33.240 ;
        RECT 4.895 33.220 5.355 33.240 ;
        RECT 5.685 33.220 6.145 33.240 ;
        RECT 6.475 33.220 6.935 33.240 ;
        RECT 7.265 33.220 7.725 33.240 ;
        RECT 8.055 33.220 8.515 33.240 ;
        RECT 8.845 33.220 9.305 33.240 ;
        RECT 9.635 33.220 10.095 33.240 ;
        RECT 10.425 33.220 10.885 33.240 ;
        RECT 11.215 33.220 11.675 33.240 ;
        RECT 12.005 33.220 12.465 33.240 ;
        RECT 12.795 33.220 13.255 33.240 ;
        RECT 13.585 33.220 14.045 33.240 ;
        RECT 14.375 33.220 14.835 33.240 ;
        RECT 15.165 33.220 15.625 33.240 ;
        RECT 15.955 33.220 16.415 33.240 ;
        RECT 16.745 33.220 17.205 33.240 ;
        RECT 17.535 33.220 17.995 33.240 ;
        RECT 18.325 33.220 18.785 33.240 ;
        RECT 2.525 33.035 18.825 33.220 ;
        RECT 2.525 33.010 3.775 33.035 ;
        RECT 4.105 33.010 4.565 33.035 ;
        RECT 4.895 33.010 5.355 33.035 ;
        RECT 5.685 33.010 6.145 33.035 ;
        RECT 6.475 33.010 6.935 33.035 ;
        RECT 7.265 33.010 7.725 33.035 ;
        RECT 8.055 33.010 8.515 33.035 ;
        RECT 8.845 33.010 9.305 33.035 ;
        RECT 9.635 33.010 10.095 33.035 ;
        RECT 10.425 33.010 10.885 33.035 ;
        RECT 11.215 33.010 11.675 33.035 ;
        RECT 12.005 33.010 12.465 33.035 ;
        RECT 12.795 33.010 13.255 33.035 ;
        RECT 13.585 33.010 14.045 33.035 ;
        RECT 14.375 33.010 14.835 33.035 ;
        RECT 15.165 33.010 15.625 33.035 ;
        RECT 15.955 33.010 16.415 33.035 ;
        RECT 16.745 33.010 17.205 33.035 ;
        RECT 17.535 33.010 17.995 33.035 ;
        RECT 18.325 33.010 18.785 33.035 ;
        RECT 2.525 31.600 2.760 33.010 ;
        RECT 3.020 32.195 3.280 32.865 ;
        RECT 3.035 31.805 3.265 32.195 ;
        RECT 3.460 31.600 3.620 33.010 ;
        RECT 3.825 32.425 4.055 32.805 ;
        RECT 3.810 31.755 4.070 32.425 ;
        RECT 4.250 31.600 4.410 33.010 ;
        RECT 4.600 32.195 4.860 32.865 ;
        RECT 4.615 31.805 4.845 32.195 ;
        RECT 5.040 31.600 5.200 33.010 ;
        RECT 5.405 32.425 5.635 32.805 ;
        RECT 5.390 31.755 5.650 32.425 ;
        RECT 5.830 31.600 5.990 33.010 ;
        RECT 6.180 32.195 6.440 32.865 ;
        RECT 6.195 31.805 6.425 32.195 ;
        RECT 6.620 31.600 6.780 33.010 ;
        RECT 6.985 32.425 7.215 32.805 ;
        RECT 6.970 31.755 7.230 32.425 ;
        RECT 7.410 31.600 7.570 33.010 ;
        RECT 7.760 32.195 8.020 32.865 ;
        RECT 7.775 31.805 8.005 32.195 ;
        RECT 8.200 31.600 8.360 33.010 ;
        RECT 8.565 32.425 8.795 32.805 ;
        RECT 8.550 31.755 8.810 32.425 ;
        RECT 8.990 31.600 9.150 33.010 ;
        RECT 9.340 32.195 9.600 32.865 ;
        RECT 9.355 31.805 9.585 32.195 ;
        RECT 9.780 31.600 9.940 33.010 ;
        RECT 10.145 32.425 10.375 32.805 ;
        RECT 10.130 31.755 10.390 32.425 ;
        RECT 10.570 31.600 10.730 33.010 ;
        RECT 10.920 32.195 11.180 32.865 ;
        RECT 10.935 31.805 11.165 32.195 ;
        RECT 11.360 31.600 11.520 33.010 ;
        RECT 11.725 32.425 11.955 32.805 ;
        RECT 11.710 31.755 11.970 32.425 ;
        RECT 12.150 31.600 12.310 33.010 ;
        RECT 12.500 32.195 12.760 32.865 ;
        RECT 12.515 31.805 12.745 32.195 ;
        RECT 12.940 31.600 13.100 33.010 ;
        RECT 13.305 32.425 13.535 32.805 ;
        RECT 13.290 31.755 13.550 32.425 ;
        RECT 13.730 31.600 13.890 33.010 ;
        RECT 14.080 32.195 14.340 32.865 ;
        RECT 14.095 31.805 14.325 32.195 ;
        RECT 14.520 31.600 14.680 33.010 ;
        RECT 14.885 32.425 15.115 32.805 ;
        RECT 14.870 31.755 15.130 32.425 ;
        RECT 15.310 31.600 15.470 33.010 ;
        RECT 15.660 32.195 15.920 32.865 ;
        RECT 15.675 31.805 15.905 32.195 ;
        RECT 16.100 31.600 16.260 33.010 ;
        RECT 16.465 32.425 16.695 32.805 ;
        RECT 16.450 31.755 16.710 32.425 ;
        RECT 16.890 31.600 17.050 33.010 ;
        RECT 17.240 32.195 17.500 32.865 ;
        RECT 17.255 31.805 17.485 32.195 ;
        RECT 17.680 31.600 17.840 33.010 ;
        RECT 18.045 32.425 18.275 32.805 ;
        RECT 18.030 31.755 18.290 32.425 ;
        RECT 18.470 31.600 18.630 33.010 ;
        RECT 18.820 32.195 19.080 32.865 ;
        RECT 18.835 31.805 19.065 32.195 ;
        RECT 2.525 31.580 3.775 31.600 ;
        RECT 4.105 31.580 4.565 31.600 ;
        RECT 4.895 31.580 5.355 31.600 ;
        RECT 5.685 31.580 6.145 31.600 ;
        RECT 6.475 31.580 6.935 31.600 ;
        RECT 7.265 31.580 7.725 31.600 ;
        RECT 8.055 31.580 8.515 31.600 ;
        RECT 8.845 31.580 9.305 31.600 ;
        RECT 9.635 31.580 10.095 31.600 ;
        RECT 10.425 31.580 10.885 31.600 ;
        RECT 11.215 31.580 11.675 31.600 ;
        RECT 12.005 31.580 12.465 31.600 ;
        RECT 12.795 31.580 13.255 31.600 ;
        RECT 13.585 31.580 14.045 31.600 ;
        RECT 14.375 31.580 14.835 31.600 ;
        RECT 15.165 31.580 15.625 31.600 ;
        RECT 15.955 31.580 16.415 31.600 ;
        RECT 16.745 31.580 17.205 31.600 ;
        RECT 17.535 31.580 17.995 31.600 ;
        RECT 18.325 31.580 18.785 31.600 ;
        RECT 2.525 31.395 18.785 31.580 ;
        RECT 2.525 31.370 3.775 31.395 ;
        RECT 4.105 31.370 4.565 31.395 ;
        RECT 4.895 31.370 5.355 31.395 ;
        RECT 5.685 31.370 6.145 31.395 ;
        RECT 6.475 31.370 6.935 31.395 ;
        RECT 7.265 31.370 7.725 31.395 ;
        RECT 8.055 31.370 8.515 31.395 ;
        RECT 8.845 31.370 9.305 31.395 ;
        RECT 9.635 31.370 10.095 31.395 ;
        RECT 10.425 31.370 10.885 31.395 ;
        RECT 11.215 31.370 11.675 31.395 ;
        RECT 12.005 31.370 12.465 31.395 ;
        RECT 12.795 31.370 13.255 31.395 ;
        RECT 13.585 31.370 14.045 31.395 ;
        RECT 14.375 31.370 14.835 31.395 ;
        RECT 15.165 31.370 15.625 31.395 ;
        RECT 15.955 31.370 16.415 31.395 ;
        RECT 16.745 31.370 17.205 31.395 ;
        RECT 17.535 31.370 17.995 31.395 ;
        RECT 18.325 31.370 18.785 31.395 ;
        RECT 2.525 31.060 2.760 31.370 ;
        RECT 3.460 31.060 3.620 31.370 ;
        RECT 4.250 31.060 4.410 31.370 ;
        RECT 5.040 31.060 5.200 31.370 ;
        RECT 5.830 31.060 5.990 31.370 ;
        RECT 6.620 31.060 6.780 31.370 ;
        RECT 7.410 31.060 7.570 31.370 ;
        RECT 8.200 31.060 8.360 31.370 ;
        RECT 8.990 31.060 9.150 31.370 ;
        RECT 9.780 31.060 9.940 31.370 ;
        RECT 10.570 31.060 10.730 31.370 ;
        RECT 11.360 31.060 11.520 31.370 ;
        RECT 12.150 31.060 12.310 31.370 ;
        RECT 12.940 31.060 13.100 31.370 ;
        RECT 13.730 31.060 13.890 31.370 ;
        RECT 14.520 31.060 14.680 31.370 ;
        RECT 15.310 31.060 15.470 31.370 ;
        RECT 16.100 31.060 16.260 31.370 ;
        RECT 16.890 31.060 17.050 31.370 ;
        RECT 17.680 31.060 17.840 31.370 ;
        RECT 18.470 31.060 18.630 31.370 ;
        RECT 2.525 31.040 3.775 31.060 ;
        RECT 4.105 31.040 4.565 31.060 ;
        RECT 4.895 31.040 5.355 31.060 ;
        RECT 5.685 31.040 6.145 31.060 ;
        RECT 6.475 31.040 6.935 31.060 ;
        RECT 7.265 31.040 7.725 31.060 ;
        RECT 8.055 31.040 8.515 31.060 ;
        RECT 8.845 31.040 9.305 31.060 ;
        RECT 9.635 31.040 10.095 31.060 ;
        RECT 10.425 31.040 10.885 31.060 ;
        RECT 11.215 31.040 11.675 31.060 ;
        RECT 12.005 31.040 12.465 31.060 ;
        RECT 12.795 31.040 13.255 31.060 ;
        RECT 13.585 31.040 14.045 31.060 ;
        RECT 14.375 31.040 14.835 31.060 ;
        RECT 15.165 31.040 15.625 31.060 ;
        RECT 15.955 31.040 16.415 31.060 ;
        RECT 16.745 31.040 17.205 31.060 ;
        RECT 17.535 31.040 17.995 31.060 ;
        RECT 18.325 31.040 18.785 31.060 ;
        RECT 2.525 30.855 18.825 31.040 ;
        RECT 2.525 30.830 3.775 30.855 ;
        RECT 4.105 30.830 4.565 30.855 ;
        RECT 4.895 30.830 5.355 30.855 ;
        RECT 5.685 30.830 6.145 30.855 ;
        RECT 6.475 30.830 6.935 30.855 ;
        RECT 7.265 30.830 7.725 30.855 ;
        RECT 8.055 30.830 8.515 30.855 ;
        RECT 8.845 30.830 9.305 30.855 ;
        RECT 9.635 30.830 10.095 30.855 ;
        RECT 10.425 30.830 10.885 30.855 ;
        RECT 11.215 30.830 11.675 30.855 ;
        RECT 12.005 30.830 12.465 30.855 ;
        RECT 12.795 30.830 13.255 30.855 ;
        RECT 13.585 30.830 14.045 30.855 ;
        RECT 14.375 30.830 14.835 30.855 ;
        RECT 15.165 30.830 15.625 30.855 ;
        RECT 15.955 30.830 16.415 30.855 ;
        RECT 16.745 30.830 17.205 30.855 ;
        RECT 17.535 30.830 17.995 30.855 ;
        RECT 18.325 30.830 18.785 30.855 ;
        RECT 2.525 29.420 2.760 30.830 ;
        RECT 3.020 30.015 3.280 30.685 ;
        RECT 3.035 29.625 3.265 30.015 ;
        RECT 3.460 29.420 3.620 30.830 ;
        RECT 3.825 30.245 4.055 30.625 ;
        RECT 3.810 29.575 4.070 30.245 ;
        RECT 4.250 29.420 4.410 30.830 ;
        RECT 4.600 30.015 4.860 30.685 ;
        RECT 4.615 29.625 4.845 30.015 ;
        RECT 5.040 29.420 5.200 30.830 ;
        RECT 5.405 30.245 5.635 30.625 ;
        RECT 5.390 29.575 5.650 30.245 ;
        RECT 5.830 29.420 5.990 30.830 ;
        RECT 6.180 30.015 6.440 30.685 ;
        RECT 6.195 29.625 6.425 30.015 ;
        RECT 6.620 29.420 6.780 30.830 ;
        RECT 6.985 30.245 7.215 30.625 ;
        RECT 6.970 29.575 7.230 30.245 ;
        RECT 7.410 29.420 7.570 30.830 ;
        RECT 7.760 30.015 8.020 30.685 ;
        RECT 7.775 29.625 8.005 30.015 ;
        RECT 8.200 29.420 8.360 30.830 ;
        RECT 8.565 30.245 8.795 30.625 ;
        RECT 8.550 29.575 8.810 30.245 ;
        RECT 8.990 29.420 9.150 30.830 ;
        RECT 9.340 30.015 9.600 30.685 ;
        RECT 9.355 29.625 9.585 30.015 ;
        RECT 9.780 29.420 9.940 30.830 ;
        RECT 10.145 30.245 10.375 30.625 ;
        RECT 10.130 29.575 10.390 30.245 ;
        RECT 10.570 29.420 10.730 30.830 ;
        RECT 10.920 30.015 11.180 30.685 ;
        RECT 10.935 29.625 11.165 30.015 ;
        RECT 11.360 29.420 11.520 30.830 ;
        RECT 11.725 30.245 11.955 30.625 ;
        RECT 11.710 29.575 11.970 30.245 ;
        RECT 12.150 29.420 12.310 30.830 ;
        RECT 12.500 30.015 12.760 30.685 ;
        RECT 12.515 29.625 12.745 30.015 ;
        RECT 12.940 29.420 13.100 30.830 ;
        RECT 13.305 30.245 13.535 30.625 ;
        RECT 13.290 29.575 13.550 30.245 ;
        RECT 13.730 29.420 13.890 30.830 ;
        RECT 14.080 30.015 14.340 30.685 ;
        RECT 14.095 29.625 14.325 30.015 ;
        RECT 14.520 29.420 14.680 30.830 ;
        RECT 14.885 30.245 15.115 30.625 ;
        RECT 14.870 29.575 15.130 30.245 ;
        RECT 15.310 29.420 15.470 30.830 ;
        RECT 15.660 30.015 15.920 30.685 ;
        RECT 15.675 29.625 15.905 30.015 ;
        RECT 16.100 29.420 16.260 30.830 ;
        RECT 16.465 30.245 16.695 30.625 ;
        RECT 16.450 29.575 16.710 30.245 ;
        RECT 16.890 29.420 17.050 30.830 ;
        RECT 17.240 30.015 17.500 30.685 ;
        RECT 17.255 29.625 17.485 30.015 ;
        RECT 17.680 29.420 17.840 30.830 ;
        RECT 18.045 30.245 18.275 30.625 ;
        RECT 18.030 29.575 18.290 30.245 ;
        RECT 18.470 29.420 18.630 30.830 ;
        RECT 18.820 30.015 19.080 30.685 ;
        RECT 18.835 29.625 19.065 30.015 ;
        RECT 2.525 29.400 3.775 29.420 ;
        RECT 4.105 29.400 4.565 29.420 ;
        RECT 4.895 29.400 5.355 29.420 ;
        RECT 5.685 29.400 6.145 29.420 ;
        RECT 6.475 29.400 6.935 29.420 ;
        RECT 7.265 29.400 7.725 29.420 ;
        RECT 8.055 29.400 8.515 29.420 ;
        RECT 8.845 29.400 9.305 29.420 ;
        RECT 9.635 29.400 10.095 29.420 ;
        RECT 10.425 29.400 10.885 29.420 ;
        RECT 11.215 29.400 11.675 29.420 ;
        RECT 12.005 29.400 12.465 29.420 ;
        RECT 12.795 29.400 13.255 29.420 ;
        RECT 13.585 29.400 14.045 29.420 ;
        RECT 14.375 29.400 14.835 29.420 ;
        RECT 15.165 29.400 15.625 29.420 ;
        RECT 15.955 29.400 16.415 29.420 ;
        RECT 16.745 29.400 17.205 29.420 ;
        RECT 17.535 29.400 17.995 29.420 ;
        RECT 18.325 29.400 18.785 29.420 ;
        RECT 2.525 29.215 18.785 29.400 ;
        RECT 2.525 29.190 3.775 29.215 ;
        RECT 4.105 29.190 4.565 29.215 ;
        RECT 4.895 29.190 5.355 29.215 ;
        RECT 5.685 29.190 6.145 29.215 ;
        RECT 6.475 29.190 6.935 29.215 ;
        RECT 7.265 29.190 7.725 29.215 ;
        RECT 8.055 29.190 8.515 29.215 ;
        RECT 8.845 29.190 9.305 29.215 ;
        RECT 9.635 29.190 10.095 29.215 ;
        RECT 10.425 29.190 10.885 29.215 ;
        RECT 11.215 29.190 11.675 29.215 ;
        RECT 12.005 29.190 12.465 29.215 ;
        RECT 12.795 29.190 13.255 29.215 ;
        RECT 13.585 29.190 14.045 29.215 ;
        RECT 14.375 29.190 14.835 29.215 ;
        RECT 15.165 29.190 15.625 29.215 ;
        RECT 15.955 29.190 16.415 29.215 ;
        RECT 16.745 29.190 17.205 29.215 ;
        RECT 17.535 29.190 17.995 29.215 ;
        RECT 18.325 29.190 18.785 29.215 ;
        RECT 2.525 28.880 2.760 29.190 ;
        RECT 3.460 28.880 3.620 29.190 ;
        RECT 4.250 28.880 4.410 29.190 ;
        RECT 5.040 28.880 5.200 29.190 ;
        RECT 5.830 28.880 5.990 29.190 ;
        RECT 6.620 28.880 6.780 29.190 ;
        RECT 7.410 28.880 7.570 29.190 ;
        RECT 8.200 28.880 8.360 29.190 ;
        RECT 8.990 28.880 9.150 29.190 ;
        RECT 9.780 28.880 9.940 29.190 ;
        RECT 10.570 28.880 10.730 29.190 ;
        RECT 11.360 28.880 11.520 29.190 ;
        RECT 12.150 28.880 12.310 29.190 ;
        RECT 12.940 28.880 13.100 29.190 ;
        RECT 13.730 28.880 13.890 29.190 ;
        RECT 14.520 28.880 14.680 29.190 ;
        RECT 15.310 28.880 15.470 29.190 ;
        RECT 16.100 28.880 16.260 29.190 ;
        RECT 16.890 28.880 17.050 29.190 ;
        RECT 17.680 28.880 17.840 29.190 ;
        RECT 18.470 28.880 18.630 29.190 ;
        RECT 2.525 28.860 3.775 28.880 ;
        RECT 4.105 28.860 4.565 28.880 ;
        RECT 4.895 28.860 5.355 28.880 ;
        RECT 5.685 28.860 6.145 28.880 ;
        RECT 6.475 28.860 6.935 28.880 ;
        RECT 7.265 28.860 7.725 28.880 ;
        RECT 8.055 28.860 8.515 28.880 ;
        RECT 8.845 28.860 9.305 28.880 ;
        RECT 9.635 28.860 10.095 28.880 ;
        RECT 10.425 28.860 10.885 28.880 ;
        RECT 11.215 28.860 11.675 28.880 ;
        RECT 12.005 28.860 12.465 28.880 ;
        RECT 12.795 28.860 13.255 28.880 ;
        RECT 13.585 28.860 14.045 28.880 ;
        RECT 14.375 28.860 14.835 28.880 ;
        RECT 15.165 28.860 15.625 28.880 ;
        RECT 15.955 28.860 16.415 28.880 ;
        RECT 16.745 28.860 17.205 28.880 ;
        RECT 17.535 28.860 17.995 28.880 ;
        RECT 18.325 28.860 18.785 28.880 ;
        RECT 2.525 28.675 18.825 28.860 ;
        RECT 2.525 28.650 3.775 28.675 ;
        RECT 4.105 28.650 4.565 28.675 ;
        RECT 4.895 28.650 5.355 28.675 ;
        RECT 5.685 28.650 6.145 28.675 ;
        RECT 6.475 28.650 6.935 28.675 ;
        RECT 7.265 28.650 7.725 28.675 ;
        RECT 8.055 28.650 8.515 28.675 ;
        RECT 8.845 28.650 9.305 28.675 ;
        RECT 9.635 28.650 10.095 28.675 ;
        RECT 10.425 28.650 10.885 28.675 ;
        RECT 11.215 28.650 11.675 28.675 ;
        RECT 12.005 28.650 12.465 28.675 ;
        RECT 12.795 28.650 13.255 28.675 ;
        RECT 13.585 28.650 14.045 28.675 ;
        RECT 14.375 28.650 14.835 28.675 ;
        RECT 15.165 28.650 15.625 28.675 ;
        RECT 15.955 28.650 16.415 28.675 ;
        RECT 16.745 28.650 17.205 28.675 ;
        RECT 17.535 28.650 17.995 28.675 ;
        RECT 18.325 28.650 18.785 28.675 ;
        RECT 2.525 27.240 2.760 28.650 ;
        RECT 3.020 27.835 3.280 28.505 ;
        RECT 3.035 27.445 3.265 27.835 ;
        RECT 3.460 27.240 3.620 28.650 ;
        RECT 3.825 28.065 4.055 28.445 ;
        RECT 3.810 27.395 4.070 28.065 ;
        RECT 4.250 27.240 4.410 28.650 ;
        RECT 4.600 27.835 4.860 28.505 ;
        RECT 4.615 27.445 4.845 27.835 ;
        RECT 5.040 27.240 5.200 28.650 ;
        RECT 5.405 28.065 5.635 28.445 ;
        RECT 5.390 27.395 5.650 28.065 ;
        RECT 5.830 27.240 5.990 28.650 ;
        RECT 6.180 27.835 6.440 28.505 ;
        RECT 6.195 27.445 6.425 27.835 ;
        RECT 6.620 27.240 6.780 28.650 ;
        RECT 6.985 28.065 7.215 28.445 ;
        RECT 6.970 27.395 7.230 28.065 ;
        RECT 7.410 27.240 7.570 28.650 ;
        RECT 7.760 27.835 8.020 28.505 ;
        RECT 7.775 27.445 8.005 27.835 ;
        RECT 8.200 27.240 8.360 28.650 ;
        RECT 8.565 28.065 8.795 28.445 ;
        RECT 8.550 27.395 8.810 28.065 ;
        RECT 8.990 27.240 9.150 28.650 ;
        RECT 9.340 27.835 9.600 28.505 ;
        RECT 9.355 27.445 9.585 27.835 ;
        RECT 9.780 27.240 9.940 28.650 ;
        RECT 10.145 28.065 10.375 28.445 ;
        RECT 10.130 27.395 10.390 28.065 ;
        RECT 10.570 27.240 10.730 28.650 ;
        RECT 10.920 27.835 11.180 28.505 ;
        RECT 10.935 27.445 11.165 27.835 ;
        RECT 11.360 27.240 11.520 28.650 ;
        RECT 11.725 28.065 11.955 28.445 ;
        RECT 11.710 27.395 11.970 28.065 ;
        RECT 12.150 27.240 12.310 28.650 ;
        RECT 12.500 27.835 12.760 28.505 ;
        RECT 12.515 27.445 12.745 27.835 ;
        RECT 12.940 27.240 13.100 28.650 ;
        RECT 13.305 28.065 13.535 28.445 ;
        RECT 13.290 27.395 13.550 28.065 ;
        RECT 13.730 27.240 13.890 28.650 ;
        RECT 14.080 27.835 14.340 28.505 ;
        RECT 14.095 27.445 14.325 27.835 ;
        RECT 14.520 27.240 14.680 28.650 ;
        RECT 14.885 28.065 15.115 28.445 ;
        RECT 14.870 27.395 15.130 28.065 ;
        RECT 15.310 27.240 15.470 28.650 ;
        RECT 15.660 27.835 15.920 28.505 ;
        RECT 15.675 27.445 15.905 27.835 ;
        RECT 16.100 27.240 16.260 28.650 ;
        RECT 16.465 28.065 16.695 28.445 ;
        RECT 16.450 27.395 16.710 28.065 ;
        RECT 16.890 27.240 17.050 28.650 ;
        RECT 17.240 27.835 17.500 28.505 ;
        RECT 17.255 27.445 17.485 27.835 ;
        RECT 17.680 27.240 17.840 28.650 ;
        RECT 18.045 28.065 18.275 28.445 ;
        RECT 18.030 27.395 18.290 28.065 ;
        RECT 18.470 27.240 18.630 28.650 ;
        RECT 18.820 27.835 19.080 28.505 ;
        RECT 18.835 27.445 19.065 27.835 ;
        RECT 2.525 27.220 3.775 27.240 ;
        RECT 4.105 27.220 4.565 27.240 ;
        RECT 4.895 27.220 5.355 27.240 ;
        RECT 5.685 27.220 6.145 27.240 ;
        RECT 6.475 27.220 6.935 27.240 ;
        RECT 7.265 27.220 7.725 27.240 ;
        RECT 8.055 27.220 8.515 27.240 ;
        RECT 8.845 27.220 9.305 27.240 ;
        RECT 9.635 27.220 10.095 27.240 ;
        RECT 10.425 27.220 10.885 27.240 ;
        RECT 11.215 27.220 11.675 27.240 ;
        RECT 12.005 27.220 12.465 27.240 ;
        RECT 12.795 27.220 13.255 27.240 ;
        RECT 13.585 27.220 14.045 27.240 ;
        RECT 14.375 27.220 14.835 27.240 ;
        RECT 15.165 27.220 15.625 27.240 ;
        RECT 15.955 27.220 16.415 27.240 ;
        RECT 16.745 27.220 17.205 27.240 ;
        RECT 17.535 27.220 17.995 27.240 ;
        RECT 18.325 27.220 18.785 27.240 ;
        RECT 2.525 27.035 18.785 27.220 ;
        RECT 2.525 27.010 3.775 27.035 ;
        RECT 4.105 27.010 4.565 27.035 ;
        RECT 4.895 27.010 5.355 27.035 ;
        RECT 5.685 27.010 6.145 27.035 ;
        RECT 6.475 27.010 6.935 27.035 ;
        RECT 7.265 27.010 7.725 27.035 ;
        RECT 8.055 27.010 8.515 27.035 ;
        RECT 8.845 27.010 9.305 27.035 ;
        RECT 9.635 27.010 10.095 27.035 ;
        RECT 10.425 27.010 10.885 27.035 ;
        RECT 11.215 27.010 11.675 27.035 ;
        RECT 12.005 27.010 12.465 27.035 ;
        RECT 12.795 27.010 13.255 27.035 ;
        RECT 13.585 27.010 14.045 27.035 ;
        RECT 14.375 27.010 14.835 27.035 ;
        RECT 15.165 27.010 15.625 27.035 ;
        RECT 15.955 27.010 16.415 27.035 ;
        RECT 16.745 27.010 17.205 27.035 ;
        RECT 17.535 27.010 17.995 27.035 ;
        RECT 18.325 27.010 18.785 27.035 ;
        RECT 2.525 26.700 2.760 27.010 ;
        RECT 3.460 26.700 3.620 27.010 ;
        RECT 4.250 26.700 4.410 27.010 ;
        RECT 5.040 26.700 5.200 27.010 ;
        RECT 5.830 26.700 5.990 27.010 ;
        RECT 6.620 26.700 6.780 27.010 ;
        RECT 7.410 26.700 7.570 27.010 ;
        RECT 8.200 26.700 8.360 27.010 ;
        RECT 8.990 26.700 9.150 27.010 ;
        RECT 9.780 26.700 9.940 27.010 ;
        RECT 10.570 26.700 10.730 27.010 ;
        RECT 11.360 26.700 11.520 27.010 ;
        RECT 12.150 26.700 12.310 27.010 ;
        RECT 12.940 26.700 13.100 27.010 ;
        RECT 13.730 26.700 13.890 27.010 ;
        RECT 14.520 26.700 14.680 27.010 ;
        RECT 15.310 26.700 15.470 27.010 ;
        RECT 16.100 26.700 16.260 27.010 ;
        RECT 16.890 26.700 17.050 27.010 ;
        RECT 17.680 26.700 17.840 27.010 ;
        RECT 18.470 26.700 18.630 27.010 ;
        RECT 2.525 26.680 3.775 26.700 ;
        RECT 4.105 26.680 4.565 26.700 ;
        RECT 4.895 26.680 5.355 26.700 ;
        RECT 5.685 26.680 6.145 26.700 ;
        RECT 6.475 26.680 6.935 26.700 ;
        RECT 7.265 26.680 7.725 26.700 ;
        RECT 8.055 26.680 8.515 26.700 ;
        RECT 8.845 26.680 9.305 26.700 ;
        RECT 9.635 26.680 10.095 26.700 ;
        RECT 10.425 26.680 10.885 26.700 ;
        RECT 11.215 26.680 11.675 26.700 ;
        RECT 12.005 26.680 12.465 26.700 ;
        RECT 12.795 26.680 13.255 26.700 ;
        RECT 13.585 26.680 14.045 26.700 ;
        RECT 14.375 26.680 14.835 26.700 ;
        RECT 15.165 26.680 15.625 26.700 ;
        RECT 15.955 26.680 16.415 26.700 ;
        RECT 16.745 26.680 17.205 26.700 ;
        RECT 17.535 26.680 17.995 26.700 ;
        RECT 18.325 26.680 18.785 26.700 ;
        RECT 2.525 26.495 18.825 26.680 ;
        RECT 2.525 26.470 3.775 26.495 ;
        RECT 4.105 26.470 4.565 26.495 ;
        RECT 4.895 26.470 5.355 26.495 ;
        RECT 5.685 26.470 6.145 26.495 ;
        RECT 6.475 26.470 6.935 26.495 ;
        RECT 7.265 26.470 7.725 26.495 ;
        RECT 8.055 26.470 8.515 26.495 ;
        RECT 8.845 26.470 9.305 26.495 ;
        RECT 9.635 26.470 10.095 26.495 ;
        RECT 10.425 26.470 10.885 26.495 ;
        RECT 11.215 26.470 11.675 26.495 ;
        RECT 12.005 26.470 12.465 26.495 ;
        RECT 12.795 26.470 13.255 26.495 ;
        RECT 13.585 26.470 14.045 26.495 ;
        RECT 14.375 26.470 14.835 26.495 ;
        RECT 15.165 26.470 15.625 26.495 ;
        RECT 15.955 26.470 16.415 26.495 ;
        RECT 16.745 26.470 17.205 26.495 ;
        RECT 17.535 26.470 17.995 26.495 ;
        RECT 18.325 26.470 18.785 26.495 ;
        RECT 2.525 25.060 2.760 26.470 ;
        RECT 3.020 25.655 3.280 26.325 ;
        RECT 3.035 25.265 3.265 25.655 ;
        RECT 3.460 25.060 3.620 26.470 ;
        RECT 3.825 25.885 4.055 26.265 ;
        RECT 3.810 25.215 4.070 25.885 ;
        RECT 4.250 25.060 4.410 26.470 ;
        RECT 4.600 25.655 4.860 26.325 ;
        RECT 4.615 25.265 4.845 25.655 ;
        RECT 5.040 25.060 5.200 26.470 ;
        RECT 5.405 25.885 5.635 26.265 ;
        RECT 5.390 25.215 5.650 25.885 ;
        RECT 5.830 25.060 5.990 26.470 ;
        RECT 6.180 25.655 6.440 26.325 ;
        RECT 6.195 25.265 6.425 25.655 ;
        RECT 6.620 25.060 6.780 26.470 ;
        RECT 6.985 25.885 7.215 26.265 ;
        RECT 6.970 25.215 7.230 25.885 ;
        RECT 7.410 25.060 7.570 26.470 ;
        RECT 7.760 25.655 8.020 26.325 ;
        RECT 7.775 25.265 8.005 25.655 ;
        RECT 8.200 25.060 8.360 26.470 ;
        RECT 8.565 25.885 8.795 26.265 ;
        RECT 8.550 25.215 8.810 25.885 ;
        RECT 8.990 25.060 9.150 26.470 ;
        RECT 9.340 25.655 9.600 26.325 ;
        RECT 9.355 25.265 9.585 25.655 ;
        RECT 9.780 25.060 9.940 26.470 ;
        RECT 10.145 25.885 10.375 26.265 ;
        RECT 10.130 25.215 10.390 25.885 ;
        RECT 10.570 25.060 10.730 26.470 ;
        RECT 10.920 25.655 11.180 26.325 ;
        RECT 10.935 25.265 11.165 25.655 ;
        RECT 11.360 25.060 11.520 26.470 ;
        RECT 11.725 25.885 11.955 26.265 ;
        RECT 11.710 25.215 11.970 25.885 ;
        RECT 12.150 25.060 12.310 26.470 ;
        RECT 12.500 25.655 12.760 26.325 ;
        RECT 12.515 25.265 12.745 25.655 ;
        RECT 12.940 25.060 13.100 26.470 ;
        RECT 13.305 25.885 13.535 26.265 ;
        RECT 13.290 25.215 13.550 25.885 ;
        RECT 13.730 25.060 13.890 26.470 ;
        RECT 14.080 25.655 14.340 26.325 ;
        RECT 14.095 25.265 14.325 25.655 ;
        RECT 14.520 25.060 14.680 26.470 ;
        RECT 14.885 25.885 15.115 26.265 ;
        RECT 14.870 25.215 15.130 25.885 ;
        RECT 15.310 25.060 15.470 26.470 ;
        RECT 15.660 25.655 15.920 26.325 ;
        RECT 15.675 25.265 15.905 25.655 ;
        RECT 16.100 25.060 16.260 26.470 ;
        RECT 16.465 25.885 16.695 26.265 ;
        RECT 16.450 25.215 16.710 25.885 ;
        RECT 16.890 25.060 17.050 26.470 ;
        RECT 17.240 25.655 17.500 26.325 ;
        RECT 17.255 25.265 17.485 25.655 ;
        RECT 17.680 25.060 17.840 26.470 ;
        RECT 18.045 25.885 18.275 26.265 ;
        RECT 18.030 25.215 18.290 25.885 ;
        RECT 18.470 25.060 18.630 26.470 ;
        RECT 18.820 25.655 19.080 26.325 ;
        RECT 18.835 25.265 19.065 25.655 ;
        RECT 2.525 25.040 3.775 25.060 ;
        RECT 4.105 25.040 4.565 25.060 ;
        RECT 4.895 25.040 5.355 25.060 ;
        RECT 5.685 25.040 6.145 25.060 ;
        RECT 6.475 25.040 6.935 25.060 ;
        RECT 7.265 25.040 7.725 25.060 ;
        RECT 8.055 25.040 8.515 25.060 ;
        RECT 8.845 25.040 9.305 25.060 ;
        RECT 9.635 25.040 10.095 25.060 ;
        RECT 10.425 25.040 10.885 25.060 ;
        RECT 11.215 25.040 11.675 25.060 ;
        RECT 12.005 25.040 12.465 25.060 ;
        RECT 12.795 25.040 13.255 25.060 ;
        RECT 13.585 25.040 14.045 25.060 ;
        RECT 14.375 25.040 14.835 25.060 ;
        RECT 15.165 25.040 15.625 25.060 ;
        RECT 15.955 25.040 16.415 25.060 ;
        RECT 16.745 25.040 17.205 25.060 ;
        RECT 17.535 25.040 17.995 25.060 ;
        RECT 18.325 25.040 18.785 25.060 ;
        RECT 2.525 24.855 18.785 25.040 ;
        RECT 2.525 24.830 3.775 24.855 ;
        RECT 4.105 24.830 4.565 24.855 ;
        RECT 4.895 24.830 5.355 24.855 ;
        RECT 5.685 24.830 6.145 24.855 ;
        RECT 6.475 24.830 6.935 24.855 ;
        RECT 7.265 24.830 7.725 24.855 ;
        RECT 8.055 24.830 8.515 24.855 ;
        RECT 8.845 24.830 9.305 24.855 ;
        RECT 9.635 24.830 10.095 24.855 ;
        RECT 10.425 24.830 10.885 24.855 ;
        RECT 11.215 24.830 11.675 24.855 ;
        RECT 12.005 24.830 12.465 24.855 ;
        RECT 12.795 24.830 13.255 24.855 ;
        RECT 13.585 24.830 14.045 24.855 ;
        RECT 14.375 24.830 14.835 24.855 ;
        RECT 15.165 24.830 15.625 24.855 ;
        RECT 15.955 24.830 16.415 24.855 ;
        RECT 16.745 24.830 17.205 24.855 ;
        RECT 17.535 24.830 17.995 24.855 ;
        RECT 18.325 24.830 18.785 24.855 ;
        RECT 2.525 24.520 2.760 24.830 ;
        RECT 3.460 24.520 3.620 24.830 ;
        RECT 4.250 24.520 4.410 24.830 ;
        RECT 5.040 24.520 5.200 24.830 ;
        RECT 5.830 24.520 5.990 24.830 ;
        RECT 6.620 24.520 6.780 24.830 ;
        RECT 7.410 24.520 7.570 24.830 ;
        RECT 8.200 24.520 8.360 24.830 ;
        RECT 8.990 24.520 9.150 24.830 ;
        RECT 9.780 24.520 9.940 24.830 ;
        RECT 10.570 24.520 10.730 24.830 ;
        RECT 11.360 24.520 11.520 24.830 ;
        RECT 12.150 24.520 12.310 24.830 ;
        RECT 12.940 24.520 13.100 24.830 ;
        RECT 13.730 24.520 13.890 24.830 ;
        RECT 14.520 24.520 14.680 24.830 ;
        RECT 15.310 24.520 15.470 24.830 ;
        RECT 16.100 24.520 16.260 24.830 ;
        RECT 16.890 24.520 17.050 24.830 ;
        RECT 17.680 24.520 17.840 24.830 ;
        RECT 18.470 24.520 18.630 24.830 ;
        RECT 2.525 24.500 3.775 24.520 ;
        RECT 4.105 24.500 4.565 24.520 ;
        RECT 4.895 24.500 5.355 24.520 ;
        RECT 5.685 24.500 6.145 24.520 ;
        RECT 6.475 24.500 6.935 24.520 ;
        RECT 7.265 24.500 7.725 24.520 ;
        RECT 8.055 24.500 8.515 24.520 ;
        RECT 8.845 24.500 9.305 24.520 ;
        RECT 9.635 24.500 10.095 24.520 ;
        RECT 10.425 24.500 10.885 24.520 ;
        RECT 11.215 24.500 11.675 24.520 ;
        RECT 12.005 24.500 12.465 24.520 ;
        RECT 12.795 24.500 13.255 24.520 ;
        RECT 13.585 24.500 14.045 24.520 ;
        RECT 14.375 24.500 14.835 24.520 ;
        RECT 15.165 24.500 15.625 24.520 ;
        RECT 15.955 24.500 16.415 24.520 ;
        RECT 16.745 24.500 17.205 24.520 ;
        RECT 17.535 24.500 17.995 24.520 ;
        RECT 18.325 24.500 18.785 24.520 ;
        RECT 2.525 24.315 18.825 24.500 ;
        RECT 2.525 24.290 3.775 24.315 ;
        RECT 4.105 24.290 4.565 24.315 ;
        RECT 4.895 24.290 5.355 24.315 ;
        RECT 5.685 24.290 6.145 24.315 ;
        RECT 6.475 24.290 6.935 24.315 ;
        RECT 7.265 24.290 7.725 24.315 ;
        RECT 8.055 24.290 8.515 24.315 ;
        RECT 8.845 24.290 9.305 24.315 ;
        RECT 9.635 24.290 10.095 24.315 ;
        RECT 10.425 24.290 10.885 24.315 ;
        RECT 11.215 24.290 11.675 24.315 ;
        RECT 12.005 24.290 12.465 24.315 ;
        RECT 12.795 24.290 13.255 24.315 ;
        RECT 13.585 24.290 14.045 24.315 ;
        RECT 14.375 24.290 14.835 24.315 ;
        RECT 15.165 24.290 15.625 24.315 ;
        RECT 15.955 24.290 16.415 24.315 ;
        RECT 16.745 24.290 17.205 24.315 ;
        RECT 17.535 24.290 17.995 24.315 ;
        RECT 18.325 24.290 18.785 24.315 ;
        RECT 2.525 22.880 2.760 24.290 ;
        RECT 3.020 23.475 3.280 24.145 ;
        RECT 3.035 23.085 3.265 23.475 ;
        RECT 3.460 22.880 3.620 24.290 ;
        RECT 3.825 23.705 4.055 24.085 ;
        RECT 3.810 23.035 4.070 23.705 ;
        RECT 4.250 22.880 4.410 24.290 ;
        RECT 4.600 23.475 4.860 24.145 ;
        RECT 4.615 23.085 4.845 23.475 ;
        RECT 5.040 22.880 5.200 24.290 ;
        RECT 5.405 23.705 5.635 24.085 ;
        RECT 5.390 23.035 5.650 23.705 ;
        RECT 5.830 22.880 5.990 24.290 ;
        RECT 6.180 23.475 6.440 24.145 ;
        RECT 6.195 23.085 6.425 23.475 ;
        RECT 6.620 22.880 6.780 24.290 ;
        RECT 6.985 23.705 7.215 24.085 ;
        RECT 6.970 23.035 7.230 23.705 ;
        RECT 7.410 22.880 7.570 24.290 ;
        RECT 7.760 23.475 8.020 24.145 ;
        RECT 7.775 23.085 8.005 23.475 ;
        RECT 8.200 22.880 8.360 24.290 ;
        RECT 8.565 23.705 8.795 24.085 ;
        RECT 8.550 23.035 8.810 23.705 ;
        RECT 8.990 22.880 9.150 24.290 ;
        RECT 9.340 23.475 9.600 24.145 ;
        RECT 9.355 23.085 9.585 23.475 ;
        RECT 9.780 22.880 9.940 24.290 ;
        RECT 10.145 23.705 10.375 24.085 ;
        RECT 10.130 23.035 10.390 23.705 ;
        RECT 10.570 22.880 10.730 24.290 ;
        RECT 10.920 23.475 11.180 24.145 ;
        RECT 10.935 23.085 11.165 23.475 ;
        RECT 11.360 22.880 11.520 24.290 ;
        RECT 11.725 23.705 11.955 24.085 ;
        RECT 11.710 23.035 11.970 23.705 ;
        RECT 12.150 22.880 12.310 24.290 ;
        RECT 12.500 23.475 12.760 24.145 ;
        RECT 12.515 23.085 12.745 23.475 ;
        RECT 12.940 22.880 13.100 24.290 ;
        RECT 13.305 23.705 13.535 24.085 ;
        RECT 13.290 23.035 13.550 23.705 ;
        RECT 13.730 22.880 13.890 24.290 ;
        RECT 14.080 23.475 14.340 24.145 ;
        RECT 14.095 23.085 14.325 23.475 ;
        RECT 14.520 22.880 14.680 24.290 ;
        RECT 14.885 23.705 15.115 24.085 ;
        RECT 14.870 23.035 15.130 23.705 ;
        RECT 15.310 22.880 15.470 24.290 ;
        RECT 15.660 23.475 15.920 24.145 ;
        RECT 15.675 23.085 15.905 23.475 ;
        RECT 16.100 22.880 16.260 24.290 ;
        RECT 16.465 23.705 16.695 24.085 ;
        RECT 16.450 23.035 16.710 23.705 ;
        RECT 16.890 22.880 17.050 24.290 ;
        RECT 17.240 23.475 17.500 24.145 ;
        RECT 17.255 23.085 17.485 23.475 ;
        RECT 17.680 22.880 17.840 24.290 ;
        RECT 18.045 23.705 18.275 24.085 ;
        RECT 18.030 23.035 18.290 23.705 ;
        RECT 18.470 22.880 18.630 24.290 ;
        RECT 18.820 23.475 19.080 24.145 ;
        RECT 18.835 23.085 19.065 23.475 ;
        RECT 2.525 22.860 3.775 22.880 ;
        RECT 4.105 22.860 4.565 22.880 ;
        RECT 4.895 22.860 5.355 22.880 ;
        RECT 5.685 22.860 6.145 22.880 ;
        RECT 6.475 22.860 6.935 22.880 ;
        RECT 7.265 22.860 7.725 22.880 ;
        RECT 8.055 22.860 8.515 22.880 ;
        RECT 8.845 22.860 9.305 22.880 ;
        RECT 9.635 22.860 10.095 22.880 ;
        RECT 10.425 22.860 10.885 22.880 ;
        RECT 11.215 22.860 11.675 22.880 ;
        RECT 12.005 22.860 12.465 22.880 ;
        RECT 12.795 22.860 13.255 22.880 ;
        RECT 13.585 22.860 14.045 22.880 ;
        RECT 14.375 22.860 14.835 22.880 ;
        RECT 15.165 22.860 15.625 22.880 ;
        RECT 15.955 22.860 16.415 22.880 ;
        RECT 16.745 22.860 17.205 22.880 ;
        RECT 17.535 22.860 17.995 22.880 ;
        RECT 18.325 22.860 18.785 22.880 ;
        RECT 2.525 22.675 18.785 22.860 ;
        RECT 2.525 22.650 3.775 22.675 ;
        RECT 4.105 22.650 4.565 22.675 ;
        RECT 4.895 22.650 5.355 22.675 ;
        RECT 5.685 22.650 6.145 22.675 ;
        RECT 6.475 22.650 6.935 22.675 ;
        RECT 7.265 22.650 7.725 22.675 ;
        RECT 8.055 22.650 8.515 22.675 ;
        RECT 8.845 22.650 9.305 22.675 ;
        RECT 9.635 22.650 10.095 22.675 ;
        RECT 10.425 22.650 10.885 22.675 ;
        RECT 11.215 22.650 11.675 22.675 ;
        RECT 12.005 22.650 12.465 22.675 ;
        RECT 12.795 22.650 13.255 22.675 ;
        RECT 13.585 22.650 14.045 22.675 ;
        RECT 14.375 22.650 14.835 22.675 ;
        RECT 15.165 22.650 15.625 22.675 ;
        RECT 15.955 22.650 16.415 22.675 ;
        RECT 16.745 22.650 17.205 22.675 ;
        RECT 17.535 22.650 17.995 22.675 ;
        RECT 18.325 22.650 18.785 22.675 ;
        RECT 2.525 18.780 2.760 22.650 ;
        RECT 19.550 22.490 20.070 53.220 ;
        RECT 20.435 22.490 20.940 54.240 ;
        RECT 2.995 21.865 19.100 22.360 ;
        RECT 19.550 21.900 20.940 22.490 ;
        RECT 3.315 21.470 3.775 21.500 ;
        RECT 4.105 21.470 4.565 21.500 ;
        RECT 4.895 21.470 5.355 21.500 ;
        RECT 5.685 21.470 6.145 21.500 ;
        RECT 6.475 21.470 6.935 21.500 ;
        RECT 7.265 21.470 7.725 21.500 ;
        RECT 8.055 21.470 8.515 21.500 ;
        RECT 8.845 21.470 9.305 21.500 ;
        RECT 9.635 21.470 10.095 21.500 ;
        RECT 10.425 21.470 10.885 21.500 ;
        RECT 11.215 21.470 11.675 21.500 ;
        RECT 12.005 21.470 12.465 21.500 ;
        RECT 12.795 21.470 13.255 21.500 ;
        RECT 13.585 21.470 14.045 21.500 ;
        RECT 14.375 21.470 14.835 21.500 ;
        RECT 15.165 21.470 15.625 21.500 ;
        RECT 15.955 21.470 16.415 21.500 ;
        RECT 16.745 21.470 17.205 21.500 ;
        RECT 17.535 21.470 17.995 21.500 ;
        RECT 18.325 21.470 18.785 21.500 ;
        RECT 3.270 21.285 18.825 21.470 ;
        RECT 3.315 21.270 3.775 21.285 ;
        RECT 4.105 21.270 4.565 21.285 ;
        RECT 4.895 21.270 5.355 21.285 ;
        RECT 5.685 21.270 6.145 21.285 ;
        RECT 6.475 21.270 6.935 21.285 ;
        RECT 7.265 21.270 7.725 21.285 ;
        RECT 8.055 21.270 8.515 21.285 ;
        RECT 8.845 21.270 9.305 21.285 ;
        RECT 9.635 21.270 10.095 21.285 ;
        RECT 10.425 21.270 10.885 21.285 ;
        RECT 11.215 21.270 11.675 21.285 ;
        RECT 12.005 21.270 12.465 21.285 ;
        RECT 12.795 21.270 13.255 21.285 ;
        RECT 13.585 21.270 14.045 21.285 ;
        RECT 14.375 21.270 14.835 21.285 ;
        RECT 15.165 21.270 15.625 21.285 ;
        RECT 15.955 21.270 16.415 21.285 ;
        RECT 16.745 21.270 17.205 21.285 ;
        RECT 17.535 21.270 17.995 21.285 ;
        RECT 18.325 21.270 18.785 21.285 ;
        RECT 3.020 20.450 3.280 21.120 ;
        RECT 3.035 20.065 3.265 20.450 ;
        RECT 3.460 19.860 3.620 21.270 ;
        RECT 3.825 20.680 4.055 21.065 ;
        RECT 3.810 20.010 4.070 20.680 ;
        RECT 4.250 19.860 4.410 21.270 ;
        RECT 4.600 20.450 4.860 21.120 ;
        RECT 4.615 20.065 4.845 20.450 ;
        RECT 5.040 19.860 5.200 21.270 ;
        RECT 5.405 20.680 5.635 21.065 ;
        RECT 5.390 20.010 5.650 20.680 ;
        RECT 5.830 19.860 5.990 21.270 ;
        RECT 6.180 20.450 6.440 21.120 ;
        RECT 6.195 20.065 6.425 20.450 ;
        RECT 6.620 19.860 6.780 21.270 ;
        RECT 6.985 20.680 7.215 21.065 ;
        RECT 6.970 20.010 7.230 20.680 ;
        RECT 7.410 19.860 7.570 21.270 ;
        RECT 7.760 20.450 8.020 21.120 ;
        RECT 7.775 20.065 8.005 20.450 ;
        RECT 8.200 19.860 8.360 21.270 ;
        RECT 8.565 20.680 8.795 21.065 ;
        RECT 8.550 20.010 8.810 20.680 ;
        RECT 8.990 19.860 9.150 21.270 ;
        RECT 9.340 20.450 9.600 21.120 ;
        RECT 9.355 20.065 9.585 20.450 ;
        RECT 9.780 19.860 9.940 21.270 ;
        RECT 10.145 20.680 10.375 21.065 ;
        RECT 10.130 20.010 10.390 20.680 ;
        RECT 10.570 19.860 10.730 21.270 ;
        RECT 10.920 20.450 11.180 21.120 ;
        RECT 10.935 20.065 11.165 20.450 ;
        RECT 11.360 19.860 11.520 21.270 ;
        RECT 11.725 20.680 11.955 21.065 ;
        RECT 11.710 20.010 11.970 20.680 ;
        RECT 12.150 19.860 12.310 21.270 ;
        RECT 12.500 20.450 12.760 21.120 ;
        RECT 12.515 20.065 12.745 20.450 ;
        RECT 12.940 19.860 13.100 21.270 ;
        RECT 13.305 20.680 13.535 21.065 ;
        RECT 13.290 20.010 13.550 20.680 ;
        RECT 13.730 19.860 13.890 21.270 ;
        RECT 14.080 20.450 14.340 21.120 ;
        RECT 14.095 20.065 14.325 20.450 ;
        RECT 14.520 19.860 14.680 21.270 ;
        RECT 14.885 20.680 15.115 21.065 ;
        RECT 14.870 20.010 15.130 20.680 ;
        RECT 15.310 19.860 15.470 21.270 ;
        RECT 15.660 20.450 15.920 21.120 ;
        RECT 15.675 20.065 15.905 20.450 ;
        RECT 16.100 19.860 16.260 21.270 ;
        RECT 16.465 20.680 16.695 21.065 ;
        RECT 16.450 20.010 16.710 20.680 ;
        RECT 16.890 19.860 17.050 21.270 ;
        RECT 17.240 20.450 17.500 21.120 ;
        RECT 17.255 20.065 17.485 20.450 ;
        RECT 17.680 19.860 17.840 21.270 ;
        RECT 18.045 20.680 18.275 21.065 ;
        RECT 18.030 20.010 18.290 20.680 ;
        RECT 18.470 19.860 18.630 21.270 ;
        RECT 18.820 20.450 19.080 21.120 ;
        RECT 18.835 20.065 19.065 20.450 ;
        RECT 3.315 19.835 3.775 19.860 ;
        RECT 4.105 19.835 4.565 19.860 ;
        RECT 4.895 19.835 5.355 19.860 ;
        RECT 5.685 19.835 6.145 19.860 ;
        RECT 6.475 19.835 6.935 19.860 ;
        RECT 7.265 19.835 7.725 19.860 ;
        RECT 8.055 19.835 8.515 19.860 ;
        RECT 8.845 19.835 9.305 19.860 ;
        RECT 9.635 19.835 10.095 19.860 ;
        RECT 10.425 19.835 10.885 19.860 ;
        RECT 11.215 19.835 11.675 19.860 ;
        RECT 12.005 19.835 12.465 19.860 ;
        RECT 12.795 19.835 13.255 19.860 ;
        RECT 13.585 19.835 14.045 19.860 ;
        RECT 14.375 19.835 14.835 19.860 ;
        RECT 15.165 19.835 15.625 19.860 ;
        RECT 15.955 19.835 16.415 19.860 ;
        RECT 16.745 19.835 17.205 19.860 ;
        RECT 17.535 19.835 17.995 19.860 ;
        RECT 18.325 19.835 18.785 19.860 ;
        RECT 3.255 19.650 18.810 19.835 ;
        RECT 3.315 19.630 3.775 19.650 ;
        RECT 4.105 19.630 4.565 19.650 ;
        RECT 4.895 19.630 5.355 19.650 ;
        RECT 5.685 19.630 6.145 19.650 ;
        RECT 6.475 19.630 6.935 19.650 ;
        RECT 7.265 19.630 7.725 19.650 ;
        RECT 8.055 19.630 8.515 19.650 ;
        RECT 8.845 19.630 9.305 19.650 ;
        RECT 9.635 19.630 10.095 19.650 ;
        RECT 10.425 19.630 10.885 19.650 ;
        RECT 11.215 19.630 11.675 19.650 ;
        RECT 12.005 19.630 12.465 19.650 ;
        RECT 12.795 19.630 13.255 19.650 ;
        RECT 13.585 19.630 14.045 19.650 ;
        RECT 14.375 19.630 14.835 19.650 ;
        RECT 15.075 19.630 15.625 19.650 ;
        RECT 15.955 19.630 16.415 19.650 ;
        RECT 16.745 19.630 17.205 19.650 ;
        RECT 17.535 19.630 17.995 19.650 ;
        RECT 18.325 19.630 18.785 19.650 ;
        RECT 3.255 18.960 14.795 19.280 ;
        RECT 2.525 18.545 10.790 18.780 ;
        RECT 0.895 18.355 2.285 18.465 ;
        RECT 0.895 18.050 10.200 18.355 ;
        RECT 0.895 17.920 2.285 18.050 ;
        RECT 0.895 -6.075 1.415 17.920 ;
        RECT 1.750 -3.160 2.285 17.920 ;
        RECT 10.555 17.700 10.790 18.545 ;
        RECT 11.015 18.025 14.900 18.365 ;
        RECT 15.075 17.700 15.265 19.630 ;
        RECT 19.550 19.275 20.070 21.900 ;
        RECT 15.465 18.960 20.070 19.275 ;
        RECT 19.550 18.485 20.070 18.960 ;
        RECT 20.435 18.485 20.940 21.900 ;
        RECT 19.550 18.360 20.940 18.485 ;
        RECT 15.480 18.025 20.940 18.360 ;
        RECT 19.550 17.940 20.940 18.025 ;
        RECT 3.290 17.365 3.750 17.595 ;
        RECT 4.080 17.365 4.540 17.595 ;
        RECT 4.870 17.365 5.330 17.595 ;
        RECT 7.000 17.365 7.460 17.595 ;
        RECT 7.790 17.365 8.250 17.595 ;
        RECT 8.580 17.365 9.040 17.595 ;
        RECT 9.370 17.365 9.830 17.595 ;
        RECT 2.955 17.160 3.140 17.175 ;
        RECT 2.955 16.160 3.240 17.160 ;
        RECT 2.955 15.940 3.140 16.160 ;
        RECT 3.435 15.955 3.590 17.365 ;
        RECT 3.785 16.555 4.045 17.225 ;
        RECT 3.800 16.160 4.030 16.555 ;
        RECT 4.225 15.955 4.380 17.365 ;
        RECT 4.590 16.765 4.820 17.160 ;
        RECT 4.580 16.095 4.840 16.765 ;
        RECT 5.015 15.955 5.170 17.365 ;
        RECT 5.365 16.555 5.625 17.225 ;
        RECT 6.700 16.555 6.960 17.225 ;
        RECT 5.380 16.160 5.610 16.555 ;
        RECT 6.720 16.160 6.950 16.555 ;
        RECT 7.145 15.955 7.300 17.365 ;
        RECT 7.510 16.770 7.740 17.160 ;
        RECT 7.490 16.100 7.750 16.770 ;
        RECT 7.935 15.955 8.090 17.365 ;
        RECT 8.280 16.555 8.540 17.225 ;
        RECT 8.300 16.160 8.530 16.555 ;
        RECT 8.725 15.955 8.880 17.365 ;
        RECT 9.090 16.765 9.320 17.160 ;
        RECT 9.055 16.160 9.320 16.765 ;
        RECT 9.055 16.095 9.315 16.160 ;
        RECT 9.515 15.955 9.670 17.365 ;
        RECT 9.865 16.555 10.125 17.225 ;
        RECT 9.880 16.160 10.110 16.555 ;
        RECT 3.290 15.940 3.750 15.955 ;
        RECT 4.080 15.940 4.540 15.955 ;
        RECT 4.870 15.940 5.330 15.955 ;
        RECT 2.955 15.750 5.370 15.940 ;
        RECT 3.290 15.725 3.750 15.750 ;
        RECT 4.080 15.725 4.540 15.750 ;
        RECT 4.870 15.725 5.330 15.750 ;
        RECT 7.000 15.725 7.460 15.955 ;
        RECT 7.790 15.725 8.250 15.955 ;
        RECT 8.580 15.725 9.040 15.955 ;
        RECT 9.370 15.725 9.830 15.955 ;
        RECT 2.895 13.595 3.155 14.265 ;
        RECT 2.485 12.695 2.745 13.365 ;
        RECT 2.510 7.265 2.745 12.695 ;
        RECT 2.935 9.155 3.135 13.595 ;
        RECT 3.430 10.450 3.615 15.725 ;
        RECT 4.130 15.485 4.800 15.515 ;
        RECT 7.145 15.485 7.300 15.725 ;
        RECT 7.935 15.485 8.090 15.725 ;
        RECT 4.130 15.330 8.090 15.485 ;
        RECT 4.130 15.255 4.800 15.330 ;
        RECT 7.935 14.540 8.090 15.330 ;
        RECT 8.725 14.870 8.880 15.725 ;
        RECT 9.515 14.870 9.670 15.725 ;
        RECT 10.455 15.445 10.895 17.700 ;
        RECT 11.500 17.365 11.960 17.595 ;
        RECT 12.290 17.365 12.750 17.595 ;
        RECT 13.080 17.365 13.540 17.595 ;
        RECT 13.870 17.365 14.330 17.595 ;
        RECT 11.195 16.555 11.455 17.225 ;
        RECT 11.220 16.160 11.450 16.555 ;
        RECT 11.645 15.955 11.800 17.365 ;
        RECT 12.010 16.770 12.240 17.160 ;
        RECT 12.000 16.100 12.260 16.770 ;
        RECT 12.435 15.955 12.590 17.365 ;
        RECT 12.775 16.555 13.035 17.225 ;
        RECT 12.800 16.160 13.030 16.555 ;
        RECT 13.225 15.955 13.380 17.365 ;
        RECT 13.590 16.765 13.820 17.160 ;
        RECT 13.565 16.095 13.825 16.765 ;
        RECT 13.570 15.955 13.825 16.095 ;
        RECT 14.015 15.955 14.170 17.365 ;
        RECT 14.360 16.555 14.620 17.225 ;
        RECT 14.380 16.160 14.610 16.555 ;
        RECT 11.475 15.740 14.365 15.955 ;
        RECT 11.500 15.725 11.960 15.740 ;
        RECT 12.290 15.725 12.750 15.740 ;
        RECT 13.080 15.725 13.540 15.740 ;
        RECT 13.870 15.725 14.330 15.740 ;
        RECT 14.975 15.435 15.360 17.700 ;
        RECT 16.000 17.365 16.460 17.595 ;
        RECT 16.790 17.365 17.250 17.595 ;
        RECT 17.580 17.365 18.040 17.595 ;
        RECT 18.370 17.365 18.830 17.595 ;
        RECT 15.695 16.555 15.955 17.225 ;
        RECT 15.720 16.160 15.950 16.555 ;
        RECT 16.155 15.955 16.310 17.365 ;
        RECT 16.510 16.770 16.740 17.160 ;
        RECT 16.500 16.100 16.760 16.770 ;
        RECT 16.945 15.955 17.100 17.365 ;
        RECT 17.275 16.555 17.535 17.225 ;
        RECT 17.300 16.160 17.530 16.555 ;
        RECT 17.735 15.955 17.890 17.365 ;
        RECT 18.090 16.765 18.320 17.160 ;
        RECT 18.065 16.095 18.325 16.765 ;
        RECT 18.090 15.955 18.320 16.095 ;
        RECT 18.525 15.955 18.680 17.365 ;
        RECT 18.860 16.555 19.120 17.225 ;
        RECT 18.880 16.160 19.110 16.555 ;
        RECT 16.000 15.945 16.460 15.955 ;
        RECT 16.790 15.945 17.250 15.955 ;
        RECT 17.580 15.945 18.830 15.955 ;
        RECT 15.990 15.740 18.850 15.945 ;
        RECT 16.000 15.725 16.460 15.740 ;
        RECT 16.790 15.725 17.250 15.740 ;
        RECT 17.580 15.725 18.830 15.740 ;
        RECT 19.550 15.510 20.070 17.940 ;
        RECT 20.435 15.275 20.940 17.940 ;
        RECT 10.590 14.870 11.260 14.955 ;
        RECT 15.000 14.870 15.155 14.875 ;
        RECT 19.595 14.870 20.765 14.995 ;
        RECT 8.725 14.715 20.765 14.870 ;
        RECT 10.590 14.695 11.260 14.715 ;
        RECT 7.935 14.385 13.970 14.540 ;
        RECT 4.055 13.295 4.845 13.305 ;
        RECT 8.525 13.295 8.680 14.385 ;
        RECT 10.605 14.125 11.275 14.200 ;
        RECT 9.315 13.970 11.275 14.125 ;
        RECT 9.315 13.295 9.470 13.970 ;
        RECT 10.605 13.940 11.275 13.970 ;
        RECT 13.815 13.295 13.970 14.385 ;
        RECT 15.000 13.295 15.155 14.715 ;
        RECT 19.595 14.585 20.765 14.715 ;
        RECT 4.055 13.075 6.990 13.295 ;
        RECT 4.055 13.070 4.845 13.075 ;
        RECT 4.080 13.065 4.845 13.070 ;
        RECT 6.230 13.065 6.990 13.075 ;
        RECT 8.380 13.065 8.840 13.295 ;
        RECT 9.170 13.065 9.630 13.295 ;
        RECT 11.320 13.065 11.780 13.295 ;
        RECT 13.470 13.065 14.330 13.295 ;
        RECT 14.660 13.065 15.520 13.295 ;
        RECT 17.210 13.065 17.670 13.295 ;
        RECT 18.000 13.065 18.460 13.295 ;
        RECT 3.800 12.555 4.030 12.905 ;
        RECT 3.785 11.885 4.045 12.555 ;
        RECT 4.230 11.745 4.385 13.065 ;
        RECT 4.580 12.250 4.840 12.920 ;
        RECT 5.950 12.550 6.180 12.905 ;
        RECT 4.590 11.905 4.820 12.250 ;
        RECT 5.930 11.880 6.190 12.550 ;
        RECT 6.380 11.745 6.535 13.065 ;
        RECT 6.730 12.260 6.990 13.065 ;
        RECT 8.075 12.260 8.335 12.930 ;
        RECT 6.740 11.905 6.970 12.260 ;
        RECT 8.100 11.905 8.330 12.260 ;
        RECT 8.525 11.745 8.680 13.065 ;
        RECT 8.890 12.555 9.120 12.905 ;
        RECT 8.880 11.885 9.140 12.555 ;
        RECT 9.315 11.745 9.470 13.065 ;
        RECT 9.680 12.260 9.940 12.930 ;
        RECT 11.040 12.560 11.270 12.905 ;
        RECT 9.680 11.905 9.910 12.260 ;
        RECT 11.030 11.890 11.290 12.560 ;
        RECT 11.465 11.745 11.640 13.065 ;
        RECT 13.140 12.905 13.400 12.940 ;
        RECT 11.830 12.560 12.060 12.905 ;
        RECT 11.815 11.890 12.075 12.560 ;
        RECT 13.140 12.270 13.420 12.905 ;
        RECT 13.190 11.905 13.420 12.270 ;
        RECT 13.815 11.745 13.970 13.065 ;
        RECT 14.380 12.555 14.610 12.905 ;
        RECT 14.365 11.885 14.625 12.555 ;
        RECT 15.000 11.745 15.170 13.065 ;
        RECT 15.555 12.255 15.815 12.925 ;
        RECT 15.570 11.905 15.800 12.255 ;
        RECT 16.905 12.250 17.165 12.920 ;
        RECT 16.930 11.905 17.160 12.250 ;
        RECT 17.365 11.745 17.520 13.065 ;
        RECT 17.720 12.575 17.950 12.905 ;
        RECT 17.710 11.905 17.970 12.575 ;
        RECT 18.155 11.745 18.310 13.065 ;
        RECT 18.485 12.250 18.745 12.920 ;
        RECT 18.510 11.905 18.740 12.250 ;
        RECT 4.080 11.515 4.540 11.745 ;
        RECT 6.230 11.515 6.690 11.745 ;
        RECT 8.380 11.515 8.840 11.745 ;
        RECT 9.170 11.515 9.630 11.745 ;
        RECT 11.320 11.515 11.780 11.745 ;
        RECT 13.470 11.515 14.330 11.745 ;
        RECT 14.660 11.515 15.520 11.745 ;
        RECT 17.210 11.515 17.670 11.745 ;
        RECT 18.000 11.515 18.460 11.745 ;
        RECT 4.105 10.755 11.280 11.210 ;
        RECT 11.465 11.000 11.640 11.515 ;
        RECT 17.365 11.000 17.520 11.515 ;
        RECT 18.155 11.000 18.310 11.515 ;
        RECT 11.465 10.825 18.310 11.000 ;
        RECT 3.430 10.265 14.340 10.450 ;
        RECT 3.390 9.580 13.865 10.085 ;
        RECT 3.630 9.155 4.080 9.255 ;
        RECT 2.935 8.955 4.080 9.155 ;
        RECT 3.630 8.865 4.080 8.955 ;
        RECT 3.630 7.565 4.080 7.955 ;
        RECT 2.485 7.005 3.155 7.265 ;
        RECT 3.760 6.470 3.940 7.565 ;
        RECT 4.465 7.540 5.965 9.580 ;
        RECT 6.825 9.110 7.285 9.340 ;
        RECT 9.225 9.315 9.685 9.325 ;
        RECT 6.545 8.935 6.775 8.950 ;
        RECT 4.460 7.245 5.965 7.540 ;
        RECT 6.335 7.950 6.775 8.935 ;
        RECT 4.460 6.680 5.975 7.245 ;
        RECT 6.335 6.505 6.620 7.950 ;
        RECT 6.985 7.790 7.140 9.110 ;
        RECT 8.900 9.095 9.685 9.315 ;
        RECT 8.900 9.085 9.640 9.095 ;
        RECT 13.480 9.085 13.940 9.315 ;
        RECT 7.335 8.535 7.565 8.950 ;
        RECT 8.900 8.935 9.130 9.085 ;
        RECT 9.675 8.935 9.935 8.945 ;
        RECT 8.900 8.925 9.175 8.935 ;
        RECT 8.945 8.575 9.175 8.925 ;
        RECT 7.335 7.950 7.680 8.535 ;
        RECT 7.420 7.865 7.680 7.950 ;
        RECT 8.885 7.935 9.175 8.575 ;
        RECT 8.885 7.905 9.145 7.935 ;
        RECT 6.825 7.560 7.285 7.790 ;
        RECT 9.325 7.775 9.480 8.880 ;
        RECT 9.675 8.275 9.965 8.935 ;
        RECT 13.190 8.930 13.450 8.945 ;
        RECT 9.735 7.935 9.965 8.275 ;
        RECT 12.630 8.275 13.450 8.930 ;
        RECT 12.630 7.925 13.430 8.275 ;
        RECT 3.310 6.210 3.980 6.470 ;
        RECT 4.265 6.165 6.620 6.505 ;
        RECT 6.985 6.465 7.140 7.560 ;
        RECT 9.225 7.545 9.685 7.775 ;
        RECT 12.630 7.245 13.270 7.925 ;
        RECT 13.625 7.765 13.780 9.085 ;
        RECT 14.155 8.925 14.340 10.265 ;
        RECT 13.990 7.925 14.340 8.925 ;
        RECT 14.700 8.190 14.875 10.825 ;
        RECT 18.920 10.470 20.785 14.155 ;
        RECT 15.465 9.570 20.785 10.470 ;
        RECT 15.630 9.080 16.090 9.310 ;
        RECT 16.420 9.080 16.880 9.310 ;
        RECT 17.210 9.080 17.670 9.310 ;
        RECT 18.000 9.080 18.460 9.310 ;
        RECT 15.335 8.270 15.595 8.940 ;
        RECT 14.155 7.920 14.340 7.925 ;
        RECT 13.480 7.675 13.940 7.765 ;
        RECT 13.480 7.535 14.195 7.675 ;
        RECT 13.525 7.415 14.195 7.535 ;
        RECT 14.670 7.520 14.930 8.190 ;
        RECT 15.350 7.920 15.580 8.270 ;
        RECT 15.770 7.760 15.925 9.080 ;
        RECT 16.140 8.570 16.370 8.920 ;
        RECT 16.130 7.900 16.390 8.570 ;
        RECT 16.560 7.760 16.715 9.080 ;
        RECT 16.915 8.270 17.175 8.940 ;
        RECT 16.930 7.920 17.160 8.270 ;
        RECT 17.350 7.760 17.505 9.080 ;
        RECT 17.720 8.570 17.950 8.920 ;
        RECT 17.705 7.900 17.965 8.570 ;
        RECT 18.140 7.760 18.295 9.080 ;
        RECT 18.495 8.270 18.755 8.940 ;
        RECT 18.510 7.920 18.740 8.270 ;
        RECT 15.630 7.530 16.090 7.760 ;
        RECT 16.420 7.530 16.880 7.760 ;
        RECT 17.210 7.530 17.670 7.760 ;
        RECT 18.000 7.530 18.460 7.760 ;
        RECT 7.370 6.680 14.915 7.245 ;
        RECT 15.770 7.200 15.925 7.530 ;
        RECT 16.560 7.200 16.715 7.530 ;
        RECT 17.350 7.200 17.505 7.530 ;
        RECT 18.135 7.200 18.290 7.530 ;
        RECT 15.770 7.045 18.290 7.200 ;
        RECT 15.775 6.860 18.215 7.045 ;
        RECT 18.920 6.690 20.785 9.570 ;
        RECT 6.925 6.205 7.595 6.465 ;
        RECT 2.540 5.480 3.940 6.015 ;
        RECT 4.265 5.260 5.185 6.165 ;
        RECT 5.375 6.015 5.965 6.020 ;
        RECT 19.715 6.015 20.785 6.690 ;
        RECT 5.375 5.480 20.785 6.015 ;
        RECT 5.510 5.475 20.785 5.480 ;
        RECT 3.025 4.680 5.185 5.260 ;
        RECT 3.020 3.020 5.180 4.200 ;
        RECT 16.685 3.850 18.845 5.030 ;
        RECT 3.020 1.360 5.180 2.540 ;
        RECT 16.685 2.190 18.845 3.370 ;
        RECT 3.020 -0.300 5.180 0.880 ;
        RECT 16.685 0.530 18.845 1.710 ;
        RECT 3.020 -1.960 5.180 -0.780 ;
        RECT 16.685 -1.130 18.845 0.050 ;
        RECT 2.150 -4.740 2.685 -3.585 ;
        RECT 3.020 -3.620 5.180 -2.440 ;
        RECT 16.685 -2.790 18.845 -1.610 ;
        RECT 2.940 -4.150 5.120 -4.070 ;
        RECT 2.940 -4.400 5.160 -4.150 ;
        RECT 2.940 -4.500 5.120 -4.400 ;
        RECT 16.685 -4.450 18.845 -3.270 ;
        RECT 19.715 -4.740 20.785 5.475 ;
        RECT 1.915 -5.270 20.785 -4.740 ;
        RECT 0.895 -6.635 20.975 -6.075 ;
        RECT 21.390 -6.970 21.885 55.145 ;
        RECT 0.540 -7.480 21.885 -6.970 ;
      LAYER met2 ;
        RECT 1.285 53.410 19.000 53.910 ;
        RECT 1.285 52.410 1.380 53.410 ;
        RECT 2.380 53.120 19.000 53.410 ;
        RECT 2.380 52.410 2.745 53.120 ;
        RECT 19.305 52.895 20.765 53.910 ;
        RECT 1.285 51.600 2.745 52.410 ;
        RECT 2.980 52.250 20.765 52.895 ;
        RECT 2.990 51.845 3.310 52.250 ;
        RECT 3.780 51.600 4.100 52.015 ;
        RECT 4.570 51.845 4.890 52.250 ;
        RECT 5.360 51.600 5.680 52.015 ;
        RECT 6.150 51.845 6.470 52.250 ;
        RECT 6.940 51.600 7.260 52.015 ;
        RECT 7.730 51.845 8.050 52.250 ;
        RECT 8.520 51.600 8.840 52.015 ;
        RECT 9.310 51.845 9.630 52.250 ;
        RECT 10.100 51.600 10.420 52.015 ;
        RECT 10.890 51.845 11.210 52.250 ;
        RECT 11.680 51.600 12.000 52.015 ;
        RECT 12.470 51.845 12.790 52.250 ;
        RECT 13.260 51.600 13.580 52.015 ;
        RECT 14.050 51.845 14.370 52.250 ;
        RECT 14.840 51.600 15.160 52.015 ;
        RECT 15.630 51.845 15.950 52.250 ;
        RECT 16.420 51.600 16.740 52.015 ;
        RECT 17.210 51.845 17.530 52.250 ;
        RECT 18.000 51.600 18.320 52.015 ;
        RECT 18.790 51.845 19.110 52.250 ;
        RECT 1.285 50.955 19.125 51.600 ;
        RECT 1.285 49.420 2.745 50.955 ;
        RECT 19.305 50.715 20.765 52.250 ;
        RECT 2.980 50.070 20.765 50.715 ;
        RECT 2.990 49.665 3.310 50.070 ;
        RECT 3.780 49.420 4.100 49.835 ;
        RECT 4.570 49.665 4.890 50.070 ;
        RECT 5.360 49.420 5.680 49.835 ;
        RECT 6.150 49.665 6.470 50.070 ;
        RECT 6.940 49.420 7.260 49.835 ;
        RECT 7.730 49.665 8.050 50.070 ;
        RECT 8.520 49.420 8.840 49.835 ;
        RECT 9.310 49.665 9.630 50.070 ;
        RECT 10.100 49.420 10.420 49.835 ;
        RECT 10.890 49.665 11.210 50.070 ;
        RECT 11.680 49.420 12.000 49.835 ;
        RECT 12.470 49.665 12.790 50.070 ;
        RECT 13.260 49.420 13.580 49.835 ;
        RECT 14.050 49.665 14.370 50.070 ;
        RECT 14.840 49.420 15.160 49.835 ;
        RECT 15.630 49.665 15.950 50.070 ;
        RECT 16.420 49.420 16.740 49.835 ;
        RECT 17.210 49.665 17.530 50.070 ;
        RECT 18.000 49.420 18.320 49.835 ;
        RECT 18.790 49.665 19.110 50.070 ;
        RECT 1.285 48.775 19.125 49.420 ;
        RECT 1.285 47.240 2.745 48.775 ;
        RECT 19.305 48.535 20.765 50.070 ;
        RECT 2.980 47.890 20.765 48.535 ;
        RECT 2.990 47.485 3.310 47.890 ;
        RECT 3.780 47.240 4.100 47.655 ;
        RECT 4.570 47.485 4.890 47.890 ;
        RECT 5.360 47.240 5.680 47.655 ;
        RECT 6.150 47.485 6.470 47.890 ;
        RECT 6.940 47.240 7.260 47.655 ;
        RECT 7.730 47.485 8.050 47.890 ;
        RECT 8.520 47.240 8.840 47.655 ;
        RECT 9.310 47.485 9.630 47.890 ;
        RECT 10.100 47.240 10.420 47.655 ;
        RECT 10.890 47.485 11.210 47.890 ;
        RECT 11.680 47.240 12.000 47.655 ;
        RECT 12.470 47.485 12.790 47.890 ;
        RECT 13.260 47.240 13.580 47.655 ;
        RECT 14.050 47.485 14.370 47.890 ;
        RECT 14.840 47.240 15.160 47.655 ;
        RECT 15.630 47.485 15.950 47.890 ;
        RECT 16.420 47.240 16.740 47.655 ;
        RECT 17.210 47.485 17.530 47.890 ;
        RECT 18.000 47.240 18.320 47.655 ;
        RECT 18.790 47.485 19.110 47.890 ;
        RECT 1.285 46.595 19.125 47.240 ;
        RECT 1.285 45.060 2.745 46.595 ;
        RECT 19.305 46.355 20.765 47.890 ;
        RECT 2.980 45.710 20.765 46.355 ;
        RECT 2.990 45.305 3.310 45.710 ;
        RECT 3.780 45.060 4.100 45.475 ;
        RECT 4.570 45.305 4.890 45.710 ;
        RECT 5.360 45.060 5.680 45.475 ;
        RECT 6.150 45.305 6.470 45.710 ;
        RECT 6.940 45.060 7.260 45.475 ;
        RECT 7.730 45.305 8.050 45.710 ;
        RECT 8.520 45.060 8.840 45.475 ;
        RECT 9.310 45.305 9.630 45.710 ;
        RECT 10.100 45.060 10.420 45.475 ;
        RECT 10.890 45.305 11.210 45.710 ;
        RECT 11.680 45.060 12.000 45.475 ;
        RECT 12.470 45.305 12.790 45.710 ;
        RECT 13.260 45.060 13.580 45.475 ;
        RECT 14.050 45.305 14.370 45.710 ;
        RECT 14.840 45.060 15.160 45.475 ;
        RECT 15.630 45.305 15.950 45.710 ;
        RECT 16.420 45.060 16.740 45.475 ;
        RECT 17.210 45.305 17.530 45.710 ;
        RECT 18.000 45.060 18.320 45.475 ;
        RECT 18.790 45.305 19.110 45.710 ;
        RECT 1.285 44.415 19.125 45.060 ;
        RECT 1.285 42.880 2.745 44.415 ;
        RECT 19.305 44.175 20.765 45.710 ;
        RECT 2.980 43.530 20.765 44.175 ;
        RECT 2.990 43.125 3.310 43.530 ;
        RECT 3.780 42.880 4.100 43.295 ;
        RECT 4.570 43.125 4.890 43.530 ;
        RECT 5.360 42.880 5.680 43.295 ;
        RECT 6.150 43.125 6.470 43.530 ;
        RECT 6.940 42.880 7.260 43.295 ;
        RECT 7.730 43.125 8.050 43.530 ;
        RECT 8.520 42.880 8.840 43.295 ;
        RECT 9.310 43.125 9.630 43.530 ;
        RECT 10.100 42.880 10.420 43.295 ;
        RECT 10.890 43.125 11.210 43.530 ;
        RECT 11.680 42.880 12.000 43.295 ;
        RECT 12.470 43.125 12.790 43.530 ;
        RECT 13.260 42.880 13.580 43.295 ;
        RECT 14.050 43.125 14.370 43.530 ;
        RECT 14.840 42.880 15.160 43.295 ;
        RECT 15.630 43.125 15.950 43.530 ;
        RECT 16.420 42.880 16.740 43.295 ;
        RECT 17.210 43.125 17.530 43.530 ;
        RECT 18.000 42.880 18.320 43.295 ;
        RECT 18.790 43.125 19.110 43.530 ;
        RECT 1.285 42.235 19.125 42.880 ;
        RECT 1.285 40.700 2.745 42.235 ;
        RECT 19.305 41.995 20.765 43.530 ;
        RECT 2.980 41.350 20.765 41.995 ;
        RECT 2.990 40.945 3.310 41.350 ;
        RECT 3.780 40.700 4.100 41.115 ;
        RECT 4.570 40.945 4.890 41.350 ;
        RECT 5.360 40.700 5.680 41.115 ;
        RECT 6.150 40.945 6.470 41.350 ;
        RECT 6.940 40.700 7.260 41.115 ;
        RECT 7.730 40.945 8.050 41.350 ;
        RECT 8.520 40.700 8.840 41.115 ;
        RECT 9.310 40.945 9.630 41.350 ;
        RECT 10.100 40.700 10.420 41.115 ;
        RECT 10.890 40.945 11.210 41.350 ;
        RECT 11.680 40.700 12.000 41.115 ;
        RECT 12.470 40.945 12.790 41.350 ;
        RECT 13.260 40.700 13.580 41.115 ;
        RECT 14.050 40.945 14.370 41.350 ;
        RECT 14.840 40.700 15.160 41.115 ;
        RECT 15.630 40.945 15.950 41.350 ;
        RECT 16.420 40.700 16.740 41.115 ;
        RECT 17.210 40.945 17.530 41.350 ;
        RECT 18.000 40.700 18.320 41.115 ;
        RECT 18.790 40.945 19.110 41.350 ;
        RECT 1.285 40.055 19.125 40.700 ;
        RECT 1.285 38.520 2.745 40.055 ;
        RECT 19.305 39.815 20.765 41.350 ;
        RECT 2.980 39.170 20.765 39.815 ;
        RECT 2.990 38.765 3.310 39.170 ;
        RECT 3.780 38.520 4.100 38.935 ;
        RECT 4.570 38.765 4.890 39.170 ;
        RECT 5.360 38.520 5.680 38.935 ;
        RECT 6.150 38.765 6.470 39.170 ;
        RECT 6.940 38.520 7.260 38.935 ;
        RECT 7.730 38.765 8.050 39.170 ;
        RECT 8.520 38.520 8.840 38.935 ;
        RECT 9.310 38.765 9.630 39.170 ;
        RECT 10.100 38.520 10.420 38.935 ;
        RECT 10.890 38.765 11.210 39.170 ;
        RECT 11.680 38.520 12.000 38.935 ;
        RECT 12.470 38.765 12.790 39.170 ;
        RECT 13.260 38.520 13.580 38.935 ;
        RECT 14.050 38.765 14.370 39.170 ;
        RECT 14.840 38.520 15.160 38.935 ;
        RECT 15.630 38.765 15.950 39.170 ;
        RECT 16.420 38.520 16.740 38.935 ;
        RECT 17.210 38.765 17.530 39.170 ;
        RECT 18.000 38.520 18.320 38.935 ;
        RECT 18.790 38.765 19.110 39.170 ;
        RECT 1.285 37.875 19.125 38.520 ;
        RECT 1.285 36.340 2.745 37.875 ;
        RECT 19.305 37.635 20.765 39.170 ;
        RECT 2.980 36.990 20.765 37.635 ;
        RECT 2.990 36.585 3.310 36.990 ;
        RECT 3.780 36.340 4.100 36.755 ;
        RECT 4.570 36.585 4.890 36.990 ;
        RECT 5.360 36.340 5.680 36.755 ;
        RECT 6.150 36.585 6.470 36.990 ;
        RECT 6.940 36.340 7.260 36.755 ;
        RECT 7.730 36.585 8.050 36.990 ;
        RECT 8.520 36.340 8.840 36.755 ;
        RECT 9.310 36.585 9.630 36.990 ;
        RECT 10.100 36.340 10.420 36.755 ;
        RECT 10.890 36.585 11.210 36.990 ;
        RECT 11.680 36.340 12.000 36.755 ;
        RECT 12.470 36.585 12.790 36.990 ;
        RECT 13.260 36.340 13.580 36.755 ;
        RECT 14.050 36.585 14.370 36.990 ;
        RECT 14.840 36.340 15.160 36.755 ;
        RECT 15.630 36.585 15.950 36.990 ;
        RECT 16.420 36.340 16.740 36.755 ;
        RECT 17.210 36.585 17.530 36.990 ;
        RECT 18.000 36.340 18.320 36.755 ;
        RECT 18.790 36.585 19.110 36.990 ;
        RECT 1.285 35.695 19.125 36.340 ;
        RECT 1.285 34.160 2.745 35.695 ;
        RECT 19.305 35.455 20.765 36.990 ;
        RECT 2.980 34.810 20.765 35.455 ;
        RECT 2.990 34.405 3.310 34.810 ;
        RECT 3.780 34.160 4.100 34.575 ;
        RECT 4.570 34.405 4.890 34.810 ;
        RECT 5.360 34.160 5.680 34.575 ;
        RECT 6.150 34.405 6.470 34.810 ;
        RECT 6.940 34.160 7.260 34.575 ;
        RECT 7.730 34.405 8.050 34.810 ;
        RECT 8.520 34.160 8.840 34.575 ;
        RECT 9.310 34.405 9.630 34.810 ;
        RECT 10.100 34.160 10.420 34.575 ;
        RECT 10.890 34.405 11.210 34.810 ;
        RECT 11.680 34.160 12.000 34.575 ;
        RECT 12.470 34.405 12.790 34.810 ;
        RECT 13.260 34.160 13.580 34.575 ;
        RECT 14.050 34.405 14.370 34.810 ;
        RECT 14.840 34.160 15.160 34.575 ;
        RECT 15.630 34.405 15.950 34.810 ;
        RECT 16.420 34.160 16.740 34.575 ;
        RECT 17.210 34.405 17.530 34.810 ;
        RECT 18.000 34.160 18.320 34.575 ;
        RECT 18.790 34.405 19.110 34.810 ;
        RECT 1.285 33.515 19.125 34.160 ;
        RECT 1.285 31.980 2.745 33.515 ;
        RECT 19.305 33.275 20.765 34.810 ;
        RECT 2.980 32.630 20.765 33.275 ;
        RECT 2.990 32.225 3.310 32.630 ;
        RECT 3.780 31.980 4.100 32.395 ;
        RECT 4.570 32.225 4.890 32.630 ;
        RECT 5.360 31.980 5.680 32.395 ;
        RECT 6.150 32.225 6.470 32.630 ;
        RECT 6.940 31.980 7.260 32.395 ;
        RECT 7.730 32.225 8.050 32.630 ;
        RECT 8.520 31.980 8.840 32.395 ;
        RECT 9.310 32.225 9.630 32.630 ;
        RECT 10.100 31.980 10.420 32.395 ;
        RECT 10.890 32.225 11.210 32.630 ;
        RECT 11.680 31.980 12.000 32.395 ;
        RECT 12.470 32.225 12.790 32.630 ;
        RECT 13.260 31.980 13.580 32.395 ;
        RECT 14.050 32.225 14.370 32.630 ;
        RECT 14.840 31.980 15.160 32.395 ;
        RECT 15.630 32.225 15.950 32.630 ;
        RECT 16.420 31.980 16.740 32.395 ;
        RECT 17.210 32.225 17.530 32.630 ;
        RECT 18.000 31.980 18.320 32.395 ;
        RECT 18.790 32.225 19.110 32.630 ;
        RECT 1.285 31.335 19.125 31.980 ;
        RECT 1.285 29.800 2.745 31.335 ;
        RECT 19.305 31.095 20.765 32.630 ;
        RECT 2.980 30.450 20.765 31.095 ;
        RECT 2.990 30.045 3.310 30.450 ;
        RECT 3.780 29.800 4.100 30.215 ;
        RECT 4.570 30.045 4.890 30.450 ;
        RECT 5.360 29.800 5.680 30.215 ;
        RECT 6.150 30.045 6.470 30.450 ;
        RECT 6.940 29.800 7.260 30.215 ;
        RECT 7.730 30.045 8.050 30.450 ;
        RECT 8.520 29.800 8.840 30.215 ;
        RECT 9.310 30.045 9.630 30.450 ;
        RECT 10.100 29.800 10.420 30.215 ;
        RECT 10.890 30.045 11.210 30.450 ;
        RECT 11.680 29.800 12.000 30.215 ;
        RECT 12.470 30.045 12.790 30.450 ;
        RECT 13.260 29.800 13.580 30.215 ;
        RECT 14.050 30.045 14.370 30.450 ;
        RECT 14.840 29.800 15.160 30.215 ;
        RECT 15.630 30.045 15.950 30.450 ;
        RECT 16.420 29.800 16.740 30.215 ;
        RECT 17.210 30.045 17.530 30.450 ;
        RECT 18.000 29.800 18.320 30.215 ;
        RECT 18.790 30.045 19.110 30.450 ;
        RECT 1.285 29.155 19.125 29.800 ;
        RECT 1.285 27.620 2.745 29.155 ;
        RECT 19.305 28.915 20.765 30.450 ;
        RECT 2.980 28.270 20.765 28.915 ;
        RECT 2.990 27.865 3.310 28.270 ;
        RECT 3.780 27.620 4.100 28.035 ;
        RECT 4.570 27.865 4.890 28.270 ;
        RECT 5.360 27.620 5.680 28.035 ;
        RECT 6.150 27.865 6.470 28.270 ;
        RECT 6.940 27.620 7.260 28.035 ;
        RECT 7.730 27.865 8.050 28.270 ;
        RECT 8.520 27.620 8.840 28.035 ;
        RECT 9.310 27.865 9.630 28.270 ;
        RECT 10.100 27.620 10.420 28.035 ;
        RECT 10.890 27.865 11.210 28.270 ;
        RECT 11.680 27.620 12.000 28.035 ;
        RECT 12.470 27.865 12.790 28.270 ;
        RECT 13.260 27.620 13.580 28.035 ;
        RECT 14.050 27.865 14.370 28.270 ;
        RECT 14.840 27.620 15.160 28.035 ;
        RECT 15.630 27.865 15.950 28.270 ;
        RECT 16.420 27.620 16.740 28.035 ;
        RECT 17.210 27.865 17.530 28.270 ;
        RECT 18.000 27.620 18.320 28.035 ;
        RECT 18.790 27.865 19.110 28.270 ;
        RECT 1.285 26.975 19.125 27.620 ;
        RECT 1.285 25.440 2.745 26.975 ;
        RECT 19.305 26.735 20.765 28.270 ;
        RECT 2.980 26.090 20.765 26.735 ;
        RECT 2.990 25.685 3.310 26.090 ;
        RECT 3.780 25.440 4.100 25.855 ;
        RECT 4.570 25.685 4.890 26.090 ;
        RECT 5.360 25.440 5.680 25.855 ;
        RECT 6.150 25.685 6.470 26.090 ;
        RECT 6.940 25.440 7.260 25.855 ;
        RECT 7.730 25.685 8.050 26.090 ;
        RECT 8.520 25.440 8.840 25.855 ;
        RECT 9.310 25.685 9.630 26.090 ;
        RECT 10.100 25.440 10.420 25.855 ;
        RECT 10.890 25.685 11.210 26.090 ;
        RECT 11.680 25.440 12.000 25.855 ;
        RECT 12.470 25.685 12.790 26.090 ;
        RECT 13.260 25.440 13.580 25.855 ;
        RECT 14.050 25.685 14.370 26.090 ;
        RECT 14.840 25.440 15.160 25.855 ;
        RECT 15.630 25.685 15.950 26.090 ;
        RECT 16.420 25.440 16.740 25.855 ;
        RECT 17.210 25.685 17.530 26.090 ;
        RECT 18.000 25.440 18.320 25.855 ;
        RECT 18.790 25.685 19.110 26.090 ;
        RECT 1.285 24.795 19.125 25.440 ;
        RECT 1.285 23.260 2.745 24.795 ;
        RECT 19.305 24.555 20.765 26.090 ;
        RECT 2.980 23.910 20.765 24.555 ;
        RECT 2.990 23.505 3.310 23.910 ;
        RECT 3.780 23.260 4.100 23.675 ;
        RECT 4.570 23.505 4.890 23.910 ;
        RECT 5.360 23.260 5.680 23.675 ;
        RECT 6.150 23.505 6.470 23.910 ;
        RECT 6.940 23.260 7.260 23.675 ;
        RECT 7.730 23.505 8.050 23.910 ;
        RECT 8.520 23.260 8.840 23.675 ;
        RECT 9.310 23.505 9.630 23.910 ;
        RECT 10.100 23.260 10.420 23.675 ;
        RECT 10.890 23.505 11.210 23.910 ;
        RECT 11.680 23.260 12.000 23.675 ;
        RECT 12.470 23.505 12.790 23.910 ;
        RECT 13.260 23.260 13.580 23.675 ;
        RECT 14.050 23.505 14.370 23.910 ;
        RECT 14.840 23.260 15.160 23.675 ;
        RECT 15.630 23.505 15.950 23.910 ;
        RECT 16.420 23.260 16.740 23.675 ;
        RECT 17.210 23.505 17.530 23.910 ;
        RECT 18.000 23.260 18.320 23.675 ;
        RECT 18.790 23.505 19.110 23.910 ;
        RECT 1.285 22.615 19.125 23.260 ;
        RECT 19.305 22.790 20.765 23.910 ;
        RECT 1.285 22.375 2.745 22.615 ;
        RECT 1.285 21.845 19.115 22.375 ;
        RECT 1.285 20.240 2.745 21.845 ;
        RECT 19.305 21.790 19.530 22.790 ;
        RECT 20.530 21.790 20.765 22.790 ;
        RECT 19.305 21.535 20.765 21.790 ;
        RECT 2.995 21.090 20.765 21.535 ;
        RECT 2.990 20.890 20.765 21.090 ;
        RECT 2.990 20.480 3.310 20.890 ;
        RECT 3.780 20.240 4.100 20.650 ;
        RECT 4.570 20.480 4.890 20.890 ;
        RECT 5.360 20.240 5.680 20.650 ;
        RECT 6.150 20.480 6.470 20.890 ;
        RECT 6.940 20.240 7.260 20.650 ;
        RECT 7.730 20.480 8.050 20.890 ;
        RECT 8.520 20.240 8.840 20.650 ;
        RECT 9.310 20.480 9.630 20.890 ;
        RECT 10.100 20.240 10.420 20.650 ;
        RECT 10.890 20.480 11.210 20.890 ;
        RECT 11.680 20.240 12.000 20.650 ;
        RECT 12.470 20.480 12.790 20.890 ;
        RECT 13.260 20.240 13.580 20.650 ;
        RECT 14.050 20.480 14.370 20.890 ;
        RECT 14.840 20.240 15.160 20.650 ;
        RECT 15.630 20.480 15.950 20.890 ;
        RECT 16.420 20.240 16.740 20.650 ;
        RECT 17.210 20.480 17.530 20.890 ;
        RECT 18.000 20.240 18.320 20.650 ;
        RECT 18.790 20.480 19.110 20.890 ;
        RECT 1.285 19.595 19.140 20.240 ;
        RECT 1.285 19.275 2.745 19.595 ;
        RECT 19.305 19.375 20.765 20.890 ;
        RECT 1.285 18.890 19.145 19.275 ;
        RECT 1.285 18.025 19.140 18.890 ;
        RECT 1.290 17.315 2.745 18.025 ;
        RECT 1.290 17.310 2.790 17.315 ;
        RECT 1.290 16.875 5.740 17.310 ;
        RECT 6.025 16.880 10.215 17.300 ;
        RECT 3.755 16.585 4.075 16.875 ;
        RECT 4.550 16.445 4.870 16.735 ;
        RECT 5.335 16.585 5.655 16.875 ;
        RECT 6.025 16.445 6.445 16.880 ;
        RECT 6.670 16.585 6.990 16.880 ;
        RECT 2.865 16.025 6.445 16.445 ;
        RECT 7.460 16.130 7.780 16.740 ;
        RECT 8.250 16.585 8.570 16.880 ;
        RECT 9.010 16.735 9.325 16.740 ;
        RECT 7.465 15.560 7.780 16.130 ;
        RECT 2.285 15.545 4.320 15.550 ;
        RECT 2.285 15.240 4.770 15.545 ;
        RECT 2.915 14.235 3.130 15.240 ;
        RECT 4.160 15.225 4.770 15.240 ;
        RECT 5.505 15.245 7.780 15.560 ;
        RECT 9.010 16.125 9.345 16.735 ;
        RECT 9.835 16.585 10.155 16.880 ;
        RECT 5.505 14.300 5.820 15.245 ;
        RECT 9.010 14.935 9.325 16.125 ;
        RECT 10.455 15.545 10.895 17.700 ;
        RECT 11.050 17.310 11.475 18.025 ;
        RECT 11.050 16.885 14.670 17.310 ;
        RECT 11.165 16.585 11.485 16.885 ;
        RECT 11.960 15.545 12.290 16.740 ;
        RECT 12.745 16.585 13.065 16.885 ;
        RECT 2.865 13.625 3.185 14.235 ;
        RECT 4.550 13.985 5.820 14.300 ;
        RECT 6.700 14.620 9.325 14.935 ;
        RECT 10.020 15.215 12.290 15.545 ;
        RECT 2.455 13.305 2.775 13.335 ;
        RECT 4.550 13.305 4.865 13.985 ;
        RECT 2.455 12.980 4.865 13.305 ;
        RECT 2.455 12.725 2.775 12.980 ;
        RECT 4.550 12.890 4.865 12.980 ;
        RECT 6.700 12.900 7.015 14.620 ;
        RECT 10.020 14.380 10.350 15.215 ;
        RECT 10.620 14.665 11.230 14.985 ;
        RECT 13.535 14.780 13.865 16.745 ;
        RECT 14.330 16.585 14.650 16.885 ;
        RECT 14.975 15.535 15.360 17.700 ;
        RECT 15.550 17.310 15.975 18.025 ;
        RECT 15.550 16.885 19.170 17.310 ;
        RECT 15.550 16.880 15.985 16.885 ;
        RECT 15.665 16.585 15.985 16.880 ;
        RECT 16.460 15.535 16.790 16.740 ;
        RECT 17.245 16.585 17.565 16.885 ;
        RECT 8.045 14.050 10.350 14.380 ;
        RECT 10.795 14.230 11.065 14.665 ;
        RECT 11.610 14.450 13.865 14.780 ;
        RECT 14.560 15.205 16.790 15.535 ;
        RECT 3.645 11.295 4.205 12.630 ;
        RECT 4.550 12.280 4.870 12.890 ;
        RECT 5.755 11.295 6.315 12.635 ;
        RECT 6.700 12.290 7.020 12.900 ;
        RECT 8.045 12.280 8.375 14.050 ;
        RECT 10.635 13.910 11.245 14.230 ;
        RECT 11.610 13.710 11.940 14.450 ;
        RECT 9.650 13.380 11.940 13.710 ;
        RECT 8.710 12.065 9.270 12.630 ;
        RECT 9.650 12.270 9.980 13.380 ;
        RECT 14.560 13.160 14.890 15.205 ;
        RECT 18.035 14.735 18.365 16.745 ;
        RECT 18.830 16.585 19.150 16.885 ;
        RECT 13.105 12.830 14.890 13.160 ;
        RECT 15.525 14.405 18.365 14.735 ;
        RECT 11.000 12.065 11.320 12.530 ;
        RECT 8.710 11.615 11.320 12.065 ;
        RECT 11.715 11.295 12.230 12.570 ;
        RECT 13.105 12.310 13.435 12.830 ;
        RECT 13.110 12.300 13.430 12.310 ;
        RECT 14.225 12.065 14.785 12.635 ;
        RECT 15.525 12.300 15.855 14.405 ;
        RECT 16.190 12.890 18.740 13.235 ;
        RECT 16.190 12.785 18.775 12.890 ;
        RECT 15.525 12.285 15.845 12.300 ;
        RECT 16.190 12.065 16.640 12.785 ;
        RECT 16.875 12.280 17.195 12.785 ;
        RECT 14.225 11.615 16.640 12.065 ;
        RECT 17.570 11.295 18.085 12.565 ;
        RECT 18.455 12.280 18.775 12.785 ;
        RECT 1.295 10.875 19.160 11.295 ;
        RECT 1.295 9.875 1.415 10.875 ;
        RECT 2.415 9.875 19.160 10.875 ;
        RECT 1.295 8.705 19.160 9.875 ;
        RECT 7.390 8.115 7.710 8.505 ;
        RECT 8.855 8.115 9.175 8.545 ;
        RECT 9.645 8.305 9.965 8.705 ;
        RECT 13.160 8.305 13.480 8.705 ;
        RECT 15.305 8.300 15.625 8.705 ;
        RECT 14.640 8.115 14.960 8.160 ;
        RECT 16.100 8.115 16.420 8.540 ;
        RECT 16.885 8.300 17.205 8.705 ;
        RECT 17.675 8.115 17.995 8.540 ;
        RECT 18.465 8.300 18.785 8.705 ;
        RECT 19.595 8.115 20.765 19.375 ;
        RECT 6.455 7.550 15.000 8.115 ;
        RECT 15.390 7.550 20.765 8.115 ;
        RECT 13.555 7.385 14.165 7.550 ;
        RECT 2.515 7.225 3.125 7.295 ;
        RECT 2.515 7.005 18.245 7.225 ;
        RECT 2.515 6.975 3.125 7.005 ;
        RECT 15.740 6.905 18.240 7.005 ;
        RECT 3.340 6.415 3.950 6.500 ;
        RECT 6.955 6.415 7.565 6.495 ;
        RECT 2.305 6.235 7.575 6.415 ;
        RECT 3.340 6.180 3.950 6.235 ;
        RECT 6.955 6.175 7.565 6.235 ;
        RECT 19.715 6.015 20.785 6.420 ;
        RECT 1.750 -4.070 2.285 6.015 ;
        RECT 2.545 5.475 20.785 6.015 ;
        RECT 1.750 -4.490 5.120 -4.070 ;
        RECT 19.715 -4.740 20.785 5.475 ;
        RECT 1.915 -5.270 20.785 -4.740 ;
  END
END follower_amp
END LIBRARY

