VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO manual_routing
  CLASS COVER ;
  FOREIGN manual_routing ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.000 BY 1.000 ;
  OBS
      LAYER met1 ;
        RECT 1655.470 232.340 1656.470 232.585 ;
        RECT 1636.760 231.840 1685.430 232.340 ;
        RECT 1655.470 231.585 1656.470 231.840 ;
        RECT 1655.470 92.340 1656.470 92.585 ;
        RECT 1636.760 91.840 1685.430 92.340 ;
        RECT 1655.470 91.585 1656.470 91.840 ;
      LAYER met2 ;
        RECT 1665.245 238.685 1713.400 240.685 ;
        RECT 1665.245 238.565 1667.245 238.685 ;
        RECT 1616.415 236.565 1667.245 238.565 ;
        RECT 1616.415 230.790 1618.415 236.565 ;
        RECT 1665.245 233.805 1667.245 236.565 ;
        RECT 1683.400 236.165 1700.260 238.165 ;
        RECT 1683.400 233.820 1685.400 236.165 ;
        RECT 1655.470 231.585 1656.470 232.585 ;
        RECT 1634.575 199.320 1635.745 200.490 ;
        RECT 1608.410 192.510 1616.415 193.510 ;
        RECT 1608.410 166.545 1609.410 192.510 ;
        RECT 1616.440 187.410 1617.610 188.580 ;
        RECT 1674.845 166.545 1675.845 233.775 ;
        RECT 1608.410 165.545 1675.845 166.545 ;
        RECT 1665.245 98.685 1713.400 100.685 ;
        RECT 1665.245 98.565 1667.245 98.685 ;
        RECT 1616.415 96.565 1667.245 98.565 ;
        RECT 1616.415 90.790 1618.415 96.565 ;
        RECT 1665.245 93.805 1667.245 96.565 ;
        RECT 1683.400 96.165 1700.260 98.165 ;
        RECT 1683.400 93.820 1685.400 96.165 ;
        RECT 1655.470 91.585 1656.470 92.585 ;
        RECT 1634.575 59.315 1635.745 60.485 ;
        RECT 1466.980 55.000 1468.255 56.270 ;
        RECT 1566.980 55.000 1568.255 56.270 ;
        RECT 944.945 29.030 948.915 30.020 ;
        RECT 944.930 15.530 948.930 29.030 ;
        RECT 1254.980 29.025 1258.950 30.020 ;
        RECT 1254.960 15.620 1258.960 29.025 ;
        RECT 1465.610 15.620 1469.610 55.000 ;
        RECT 944.930 11.530 1074.995 15.530 ;
        RECT 1070.995 2.000 1074.995 11.530 ;
        RECT 1180.940 11.620 1258.960 15.620 ;
        RECT 1290.870 11.620 1469.610 15.620 ;
        RECT 1180.940 2.000 1184.940 11.620 ;
        RECT 1290.870 2.000 1294.870 11.620 ;
        RECT 1565.595 8.840 1569.595 55.000 ;
        RECT 1608.410 52.510 1616.415 53.510 ;
        RECT 1608.410 26.545 1609.410 52.510 ;
        RECT 1616.440 47.410 1617.610 48.580 ;
        RECT 1674.845 26.545 1675.845 93.775 ;
        RECT 1608.410 25.545 1675.845 26.545 ;
        RECT 1400.895 4.840 1569.595 8.840 ;
        RECT 1400.895 2.000 1404.895 4.840 ;
        RECT 1068.340 0.000 1077.320 2.000 ;
        RECT 1178.340 0.000 1187.320 2.000 ;
        RECT 1288.340 0.000 1297.320 2.000 ;
        RECT 1398.340 0.000 1407.320 2.000 ;
      LAYER met3 ;
        RECT 796.680 276.920 1713.400 286.920 ;
        RECT 796.680 262.630 1700.260 272.630 ;
        RECT 798.155 260.400 1609.205 261.900 ;
        RECT 798.155 210.880 799.655 260.400 ;
        RECT 1108.340 258.305 1607.140 259.805 ;
        RECT 1108.340 210.880 1109.840 258.305 ;
        RECT 798.040 208.780 800.140 210.880 ;
        RECT 1108.040 208.780 1110.140 210.880 ;
        RECT 1416.645 177.830 1418.205 178.830 ;
        RECT 1516.695 177.830 1518.255 178.830 ;
        RECT 1416.645 176.675 1417.645 177.830 ;
        RECT 1516.695 176.675 1517.695 177.830 ;
        RECT 1416.645 175.675 1418.220 176.675 ;
        RECT 1516.695 175.675 1518.270 176.675 ;
        RECT 1416.645 87.460 1418.205 88.460 ;
        RECT 1516.695 87.460 1518.255 88.460 ;
        RECT 1416.645 86.560 1417.645 87.460 ;
        RECT 1516.695 86.560 1517.695 87.460 ;
        RECT 1416.645 85.560 1418.220 86.560 ;
        RECT 1516.695 85.560 1518.270 86.560 ;
        RECT 1605.640 60.675 1607.140 258.305 ;
        RECT 1607.705 200.645 1609.205 260.400 ;
        RECT 1655.470 231.585 1656.470 232.585 ;
        RECT 1607.705 200.470 1635.145 200.645 ;
        RECT 1607.705 199.340 1635.725 200.470 ;
        RECT 1607.705 199.145 1635.145 199.340 ;
        RECT 1690.260 188.990 1700.260 262.630 ;
        RECT 1617.045 188.560 1700.260 188.990 ;
        RECT 1616.460 187.430 1700.260 188.560 ;
        RECT 1617.045 186.990 1700.260 187.430 ;
        RECT 1655.470 91.585 1656.470 92.585 ;
        RECT 1605.640 60.465 1635.155 60.675 ;
        RECT 1605.640 59.335 1635.725 60.465 ;
        RECT 1605.640 59.175 1635.155 59.335 ;
        RECT 1690.260 48.990 1700.260 186.990 ;
        RECT 1617.045 48.560 1700.260 48.990 ;
        RECT 1616.460 47.430 1700.260 48.560 ;
        RECT 1617.045 46.990 1700.260 47.430 ;
        RECT 812.120 30.750 814.900 31.745 ;
        RECT 812.120 30.110 878.405 30.750 ;
        RECT 812.120 28.965 814.900 30.110 ;
        RECT 946.555 30.000 947.315 31.295 ;
        RECT 1122.145 30.750 1124.925 31.745 ;
        RECT 1122.145 30.110 1188.430 30.750 ;
        RECT 944.965 28.070 948.895 30.000 ;
        RECT 1122.145 28.965 1124.925 30.110 ;
        RECT 1256.555 30.000 1257.315 31.295 ;
        RECT 1255.000 28.070 1258.930 30.000 ;
        RECT 1690.260 17.400 1700.260 46.990 ;
        RECT 1703.400 30.400 1713.400 276.920 ;
        RECT 1703.400 20.400 2495.655 30.400 ;
        RECT 1690.260 8.580 2365.645 17.400 ;
        RECT 1690.260 7.400 2365.655 8.580 ;
        RECT 2291.860 0.000 2315.760 7.400 ;
        RECT 2341.755 0.000 2365.655 7.400 ;
        RECT 2421.860 0.000 2445.760 20.400 ;
        RECT 2471.755 0.000 2495.655 20.400 ;
      LAYER met4 ;
        RECT 800.215 276.920 807.685 286.920 ;
        RECT 1110.215 276.920 1117.685 286.920 ;
        RECT 809.890 262.630 817.360 272.630 ;
        RECT 1119.890 262.630 1127.360 272.630 ;
        RECT 1410.190 215.850 1426.495 217.760 ;
        RECT 798.040 208.780 800.140 210.880 ;
        RECT 1108.040 208.780 1110.140 210.880 ;
        RECT 801.600 123.835 805.980 125.015 ;
        RECT 1111.560 123.835 1115.940 125.015 ;
        RECT 811.570 119.230 815.950 120.410 ;
        RECT 1121.530 119.230 1125.910 120.410 ;
        RECT 812.120 28.965 814.900 31.745 ;
        RECT 1085.460 2.150 1093.300 37.840 ;
        RECT 1122.145 28.965 1124.925 31.745 ;
        RECT 1395.460 2.150 1403.300 37.840 ;
        RECT 1410.190 11.760 1412.100 215.850 ;
        RECT 1413.895 212.450 1419.910 214.360 ;
        RECT 1413.895 2.060 1415.805 212.450 ;
        RECT 1418.000 211.255 1419.910 212.450 ;
        RECT 1424.585 211.255 1426.495 215.850 ;
        RECT 1495.850 211.255 1498.655 272.630 ;
        RECT 1499.510 211.255 1502.610 286.920 ;
        RECT 1510.190 215.850 1526.495 217.760 ;
        RECT 1510.190 11.760 1512.100 215.850 ;
        RECT 1513.895 212.450 1519.910 214.360 ;
        RECT 1513.895 2.060 1515.805 212.450 ;
        RECT 1518.000 211.255 1519.910 212.450 ;
        RECT 1524.585 211.255 1526.495 215.850 ;
        RECT 1595.850 211.255 1598.655 272.630 ;
        RECT 1599.510 211.255 1602.610 286.920 ;
        RECT 1649.430 159.560 1651.430 272.630 ;
        RECT 1652.980 159.560 1654.570 286.920 ;
        RECT 1655.345 159.560 1656.575 232.960 ;
        RECT 1652.965 11.760 1654.610 100.005 ;
        RECT 1655.345 2.060 1656.575 100.005 ;
      LAYER met5 ;
        RECT 800.215 232.235 807.685 286.920 ;
        RECT 809.890 232.235 817.360 272.630 ;
        RECT 1110.215 232.235 1117.685 286.920 ;
        RECT 1119.890 232.235 1127.360 272.630 ;
        RECT 801.480 123.625 806.100 125.225 ;
        RECT 1111.440 123.625 1116.060 125.225 ;
        RECT 811.450 119.020 816.070 120.620 ;
        RECT 1121.410 119.020 1126.030 120.620 ;
        RECT 812.000 28.845 815.020 31.865 ;
        RECT 1085.460 30.000 1093.300 37.840 ;
        RECT 1075.835 19.760 1083.675 30.000 ;
        RECT 1122.025 28.845 1125.045 31.865 ;
        RECT 1395.460 30.000 1403.300 37.840 ;
        RECT 1385.835 19.760 1393.675 30.000 ;
        RECT 798.400 11.760 1688.800 19.760 ;
        RECT 798.405 2.060 1688.800 10.060 ;
  END
END manual_routing
END LIBRARY

