`default_nettype none

module panamax_fpga_top (
    `ifdef USE_POWER_PINS
    inout wire DVPWR,    // Digital 1.8V supply
    inout wire DVGND,    // Digital ground
    inout wire AVPWR,    // Analog 3.3V supply
    inout wire AVGND,    // Analog ground
    `endif /* USE_POWER_PINS */
	
    input wire	[7:0] product_id,
    input wire	[31:0] project_id,
    
	input wire	select_tie_lo_esd,
	input wire	select_in,
	input wire	select_tie_hi_esd,
	output wire	select_enable_vddio,
	output wire	select_slow,
	inout wire	select_pad_a_esd_0_h,
	inout wire	select_pad_a_esd_1_h,
	inout wire	select_pad_a_noesd_h,
	output wire	select_analog_en,
	output wire	select_analog_pol,
	output wire	select_inp_dis,
	output wire	select_enable_inp_h,
	output wire	select_enable_h,
	output wire	select_hld_h_n,
	output wire	select_analog_sel,
	output wire	[2:0]	select_dm,
	output wire	select_hld_ovr,
	output wire	select_out,
	output wire	select_enable_vswitch_h,
	output wire	select_enable_vdda_h,
	output wire	select_vtrip_sel,
	output wire	select_ib_mode_sel,
	output wire	select_oe_n,
	input wire	select_in_h,
	input wire	select_zero,
	input wire	select_one,
	output wire	resetb_tie_weak_hi_h,
	output wire	resetb_disable_pullup_h,
	input wire	resetb_tie_hi_esd,
	input wire	resetb_xres_h_n,
	input wire	resetb_xres_n,
	input wire	resetb_tie_lo_esd,
	output wire	resetb_inp_sel_h,
	output wire	resetb_en_vddio_sig_h,
	output wire	resetb_filt_in_h,
	inout wire	resetb_pad_a_esd_h,
	output wire	resetb_pullup_h,
	output wire	resetb_enable_h,
	output wire	resetb_enable_vddio,
	input wire	gpio8_0_tie_lo_esd,
	input wire	gpio8_0_in,
	input wire	gpio8_0_tie_hi_esd,
	output wire	gpio8_0_enable_vddio,
	output wire	gpio8_0_slow,
	inout wire	gpio8_0_pad_a_esd_0_h,
	inout wire	gpio8_0_pad_a_esd_1_h,
	inout wire	gpio8_0_pad_a_noesd_h,
	output wire	gpio8_0_analog_en,
	output wire	gpio8_0_analog_pol,
	output wire	gpio8_0_inp_dis,
	output wire	gpio8_0_enable_inp_h,
	output wire	gpio8_0_enable_h,
	output wire	gpio8_0_hld_h_n,
	output wire	gpio8_0_analog_sel,
	output wire	[2:0]	gpio8_0_dm,
	output wire	gpio8_0_hld_ovr,
	output wire	gpio8_0_out,
	output wire	gpio8_0_enable_vswitch_h,
	output wire	gpio8_0_enable_vdda_h,
	output wire	gpio8_0_vtrip_sel,
	output wire	gpio8_0_ib_mode_sel,
	output wire	gpio8_0_oe_n,
	input wire	gpio8_0_in_h,
	input wire	gpio8_0_zero,
	input wire	gpio8_0_one,
	input wire	gpio8_1_tie_lo_esd,
	input wire	gpio8_1_in,
	input wire	gpio8_1_tie_hi_esd,
	output wire	gpio8_1_enable_vddio,
	output wire	gpio8_1_slow,
	inout wire	gpio8_1_pad_a_esd_0_h,
	inout wire	gpio8_1_pad_a_esd_1_h,
	inout wire	gpio8_1_pad_a_noesd_h,
	output wire	gpio8_1_analog_en,
	output wire	gpio8_1_analog_pol,
	output wire	gpio8_1_inp_dis,
	output wire	gpio8_1_enable_inp_h,
	output wire	gpio8_1_enable_h,
	output wire	gpio8_1_hld_h_n,
	output wire	gpio8_1_analog_sel,
	output wire	[2:0]	gpio8_1_dm,
	output wire	gpio8_1_hld_ovr,
	output wire	gpio8_1_out,
	output wire	gpio8_1_enable_vswitch_h,
	output wire	gpio8_1_enable_vdda_h,
	output wire	gpio8_1_vtrip_sel,
	output wire	gpio8_1_ib_mode_sel,
	output wire	gpio8_1_oe_n,
	input wire	gpio8_1_in_h,
	input wire	gpio8_1_zero,
	input wire	gpio8_1_one,
	input wire	gpio8_2_tie_lo_esd,
	input wire	gpio8_2_in,
	input wire	gpio8_2_tie_hi_esd,
	output wire	gpio8_2_enable_vddio,
	output wire	gpio8_2_slow,
	inout wire	gpio8_2_pad_a_esd_0_h,
	inout wire	gpio8_2_pad_a_esd_1_h,
	inout wire	gpio8_2_pad_a_noesd_h,
	output wire	gpio8_2_analog_en,
	output wire	gpio8_2_analog_pol,
	output wire	gpio8_2_inp_dis,
	output wire	gpio8_2_enable_inp_h,
	output wire	gpio8_2_enable_h,
	output wire	gpio8_2_hld_h_n,
	output wire	gpio8_2_analog_sel,
	output wire	[2:0]	gpio8_2_dm,
	output wire	gpio8_2_hld_ovr,
	output wire	gpio8_2_out,
	output wire	gpio8_2_enable_vswitch_h,
	output wire	gpio8_2_enable_vdda_h,
	output wire	gpio8_2_vtrip_sel,
	output wire	gpio8_2_ib_mode_sel,
	output wire	gpio8_2_oe_n,
	input wire	gpio8_2_in_h,
	input wire	gpio8_2_zero,
	input wire	gpio8_2_one,
	input wire	gpio8_3_tie_lo_esd,
	input wire	gpio8_3_in,
	input wire	gpio8_3_tie_hi_esd,
	output wire	gpio8_3_enable_vddio,
	output wire	gpio8_3_slow,
	inout wire	gpio8_3_pad_a_esd_0_h,
	inout wire	gpio8_3_pad_a_esd_1_h,
	inout wire	gpio8_3_pad_a_noesd_h,
	output wire	gpio8_3_analog_en,
	output wire	gpio8_3_analog_pol,
	output wire	gpio8_3_inp_dis,
	output wire	gpio8_3_enable_inp_h,
	output wire	gpio8_3_enable_h,
	output wire	gpio8_3_hld_h_n,
	output wire	gpio8_3_analog_sel,
	output wire	[2:0]	gpio8_3_dm,
	output wire	gpio8_3_hld_ovr,
	output wire	gpio8_3_out,
	output wire	gpio8_3_enable_vswitch_h,
	output wire	gpio8_3_enable_vdda_h,
	output wire	gpio8_3_vtrip_sel,
	output wire	gpio8_3_ib_mode_sel,
	output wire	gpio8_3_oe_n,
	input wire	gpio8_3_in_h,
	input wire	gpio8_3_zero,
	input wire	gpio8_3_one,
	inout wire	xi0_core,
	inout wire	xo0_core,
	inout wire	xi1_core,
	inout wire	xo1_core,
	input wire	gpio8_4_tie_lo_esd,
	input wire	gpio8_4_in,
	input wire	gpio8_4_tie_hi_esd,
	output wire	gpio8_4_enable_vddio,
	output wire	gpio8_4_slow,
	inout wire	gpio8_4_pad_a_esd_0_h,
	inout wire	gpio8_4_pad_a_esd_1_h,
	inout wire	gpio8_4_pad_a_noesd_h,
	output wire	gpio8_4_analog_en,
	output wire	gpio8_4_analog_pol,
	output wire	gpio8_4_inp_dis,
	output wire	gpio8_4_enable_inp_h,
	output wire	gpio8_4_enable_h,
	output wire	gpio8_4_hld_h_n,
	output wire	gpio8_4_analog_sel,
	output wire	[2:0]	gpio8_4_dm,
	output wire	gpio8_4_hld_ovr,
	output wire	gpio8_4_out,
	output wire	gpio8_4_enable_vswitch_h,
	output wire	gpio8_4_enable_vdda_h,
	output wire	gpio8_4_vtrip_sel,
	output wire	gpio8_4_ib_mode_sel,
	output wire	gpio8_4_oe_n,
	input wire	gpio8_4_in_h,
	input wire	gpio8_4_zero,
	input wire	gpio8_4_one,
	input wire	gpio8_5_tie_lo_esd,
	input wire	gpio8_5_in,
	input wire	gpio8_5_tie_hi_esd,
	output wire	gpio8_5_enable_vddio,
	output wire	gpio8_5_slow,
	inout wire	gpio8_5_pad_a_esd_0_h,
	inout wire	gpio8_5_pad_a_esd_1_h,
	inout wire	gpio8_5_pad_a_noesd_h,
	output wire	gpio8_5_analog_en,
	output wire	gpio8_5_analog_pol,
	output wire	gpio8_5_inp_dis,
	output wire	gpio8_5_enable_inp_h,
	output wire	gpio8_5_enable_h,
	output wire	gpio8_5_hld_h_n,
	output wire	gpio8_5_analog_sel,
	output wire	[2:0]	gpio8_5_dm,
	output wire	gpio8_5_hld_ovr,
	output wire	gpio8_5_out,
	output wire	gpio8_5_enable_vswitch_h,
	output wire	gpio8_5_enable_vdda_h,
	output wire	gpio8_5_vtrip_sel,
	output wire	gpio8_5_ib_mode_sel,
	output wire	gpio8_5_oe_n,
	input wire	gpio8_5_in_h,
	input wire	gpio8_5_zero,
	input wire	gpio8_5_one,
	input wire	gpio8_6_tie_lo_esd,
	input wire	gpio8_6_in,
	input wire	gpio8_6_tie_hi_esd,
	output wire	gpio8_6_enable_vddio,
	output wire	gpio8_6_slow,
	inout wire	gpio8_6_pad_a_esd_0_h,
	inout wire	gpio8_6_pad_a_esd_1_h,
	inout wire	gpio8_6_pad_a_noesd_h,
	output wire	gpio8_6_analog_en,
	output wire	gpio8_6_analog_pol,
	output wire	gpio8_6_inp_dis,
	output wire	gpio8_6_enable_inp_h,
	output wire	gpio8_6_enable_h,
	output wire	gpio8_6_hld_h_n,
	output wire	gpio8_6_analog_sel,
	output wire	[2:0]	gpio8_6_dm,
	output wire	gpio8_6_hld_ovr,
	output wire	gpio8_6_out,
	output wire	gpio8_6_enable_vswitch_h,
	output wire	gpio8_6_enable_vdda_h,
	output wire	gpio8_6_vtrip_sel,
	output wire	gpio8_6_ib_mode_sel,
	output wire	gpio8_6_oe_n,
	input wire	gpio8_6_in_h,
	input wire	gpio8_6_zero,
	input wire	gpio8_6_one,
	input wire	gpio8_7_tie_lo_esd,
	input wire	gpio8_7_in,
	input wire	gpio8_7_tie_hi_esd,
	output wire	gpio8_7_enable_vddio,
	output wire	gpio8_7_slow,
	inout wire	gpio8_7_pad_a_esd_0_h,
	inout wire	gpio8_7_pad_a_esd_1_h,
	inout wire	gpio8_7_pad_a_noesd_h,
	output wire	gpio8_7_analog_en,
	output wire	gpio8_7_analog_pol,
	output wire	gpio8_7_inp_dis,
	output wire	gpio8_7_enable_inp_h,
	output wire	gpio8_7_enable_h,
	output wire	gpio8_7_hld_h_n,
	output wire	gpio8_7_analog_sel,
	output wire	[2:0]	gpio8_7_dm,
	output wire	gpio8_7_hld_ovr,
	output wire	gpio8_7_out,
	output wire	gpio8_7_enable_vswitch_h,
	output wire	gpio8_7_enable_vdda_h,
	output wire	gpio8_7_vtrip_sel,
	output wire	gpio8_7_ib_mode_sel,
	output wire	gpio8_7_oe_n,
	input wire	gpio8_7_in_h,
	input wire	gpio8_7_zero,
	input wire	gpio8_7_one,
	input wire	pwrdet_out2_vddio_hv,
	input wire	pwrdet_out1_vddd_hv,
	output wire	pwrdet_in1_vddio_hv,
	output wire	pwrdet_in2_vddd_hv,
	output wire	pwrdet_in1_vddd_hv,
	input wire	pwrdet_out1_vddio_hv,
	input wire	pwrdet_out2_vddd_hv,
	input wire	pwrdet_out3_vddd_hv,
	input wire	pwrdet_vddio_present_vddd_hv,
	input wire	pwrdet_out3_vddio_hv,
	input wire	pwrdet_tie_lo_esd,
	output wire	pwrdet_in3_vddd_hv,
	input wire	pwrdet_vddd_present_vddio_hv,
	output wire	pwrdet_in2_vddio_hv,
	output wire	pwrdet_in3_vddio_hv,
	output wire	pwrdet_rst_por_hv_n,
	inout wire	sio_vinref_dft,
	inout wire	sio_voutref_dft,
	output wire	[1:0]	sio_vref_sel,
	output wire	sio_enable_vdda_h,
	output wire	sio_dft_refgen,
	output wire	[2:0]	sio_voh_sel,
	inout wire	amuxbus_a_n,
	inout wire	amuxbus_b_n,
	inout wire	sio_amuxbus_b,
	inout wire	sio_amuxbus_a,
	output wire	sio_vreg_en_refgen,
	output wire	sio_ibuf_sel_refgen,
	output wire	sio_vohref,
	output wire	sio_hld_h_n_refgen,
	output wire	sio_vtrip_sel_refgen,
	output wire	[1:0]	sio_pad_a_esd_0_h,
	output wire	[1:0]	sio_pad_a_noesd_h,
	output wire	[1:0]	sio_inp_dis,
	input wire	[1:0]	sio_tie_lo_esd,
	output wire	[1:0]	sio_out,
	output wire	[1:0]	sio_vtrip_sel,
	output wire	[1:0]	sio_ibuf_sel,
	output wire	[1:0]	sio_hld_h_n,
	output wire	[1:0]	sio_hld_ovr,
	input wire	[1:0]	sio_in,
	input wire	[1:0]	sio_in_h,
	output wire	[1:0]	sio_oe_n,
	output wire	[1:0]	sio_slow,
	output wire	[1:0]	sio_vreg_en,
	output wire	sio_enable_h,
	output wire	[2:0]	sio_dm1,
	inout wire	[1:0]	sio_pad_a_esd_1_h,
	output wire	[2:0]	sio_dm0,
	output wire	muxsplit_se_hld_vdda_h_n,
	output wire	muxsplit_se_enable_vdda_h,
	output wire	muxsplit_se_switch_aa_sl,
	output wire	muxsplit_se_switch_aa_s0,
	output wire	muxsplit_se_switch_bb_s0,
	output wire	muxsplit_se_switch_bb_sl,
	output wire	muxsplit_se_switch_bb_sr,
	output wire	muxsplit_se_switch_aa_sr,
	input wire	gpio0_0_tie_lo_esd,
	input wire	gpio0_0_in,
	input wire	gpio0_0_tie_hi_esd,
	output wire	gpio0_0_enable_vddio,
	output wire	gpio0_0_slow,
	inout wire	gpio0_0_pad_a_esd_0_h,
	inout wire	gpio0_0_pad_a_esd_1_h,
	inout wire	gpio0_0_pad_a_noesd_h,
	output wire	gpio0_0_analog_en,
	output wire	gpio0_0_analog_pol,
	output wire	gpio0_0_inp_dis,
	output wire	gpio0_0_enable_inp_h,
	output wire	gpio0_0_enable_h,
	output wire	gpio0_0_hld_h_n,
	output wire	gpio0_0_analog_sel,
	output wire	[2:0]	gpio0_0_dm,
	output wire	gpio0_0_hld_ovr,
	output wire	gpio0_0_out,
	output wire	gpio0_0_enable_vswitch_h,
	output wire	gpio0_0_enable_vdda_h,
	output wire	gpio0_0_vtrip_sel,
	output wire	gpio0_0_ib_mode_sel,
	output wire	gpio0_0_oe_n,
	input wire	gpio0_0_in_h,
	input wire	gpio0_0_zero,
	input wire	gpio0_0_one,
	input wire	gpio0_1_tie_lo_esd,
	input wire	gpio0_1_in,
	input wire	gpio0_1_tie_hi_esd,
	output wire	gpio0_1_enable_vddio,
	output wire	gpio0_1_slow,
	inout wire	gpio0_1_pad_a_esd_0_h,
	inout wire	gpio0_1_pad_a_esd_1_h,
	inout wire	gpio0_1_pad_a_noesd_h,
	output wire	gpio0_1_analog_en,
	output wire	gpio0_1_analog_pol,
	output wire	gpio0_1_inp_dis,
	output wire	gpio0_1_enable_inp_h,
	output wire	gpio0_1_enable_h,
	output wire	gpio0_1_hld_h_n,
	output wire	gpio0_1_analog_sel,
	output wire	[2:0]	gpio0_1_dm,
	output wire	gpio0_1_hld_ovr,
	output wire	gpio0_1_out,
	output wire	gpio0_1_enable_vswitch_h,
	output wire	gpio0_1_enable_vdda_h,
	output wire	gpio0_1_vtrip_sel,
	output wire	gpio0_1_ib_mode_sel,
	output wire	gpio0_1_oe_n,
	input wire	gpio0_1_in_h,
	input wire	gpio0_1_zero,
	input wire	gpio0_1_one,
	input wire	gpio0_2_tie_lo_esd,
	input wire	gpio0_2_in,
	input wire	gpio0_2_tie_hi_esd,
	output wire	gpio0_2_enable_vddio,
	output wire	gpio0_2_slow,
	inout wire	gpio0_2_pad_a_esd_0_h,
	inout wire	gpio0_2_pad_a_esd_1_h,
	inout wire	gpio0_2_pad_a_noesd_h,
	output wire	gpio0_2_analog_en,
	output wire	gpio0_2_analog_pol,
	output wire	gpio0_2_inp_dis,
	output wire	gpio0_2_enable_inp_h,
	output wire	gpio0_2_enable_h,
	output wire	gpio0_2_hld_h_n,
	output wire	gpio0_2_analog_sel,
	output wire	[2:0]	gpio0_2_dm,
	output wire	gpio0_2_hld_ovr,
	output wire	gpio0_2_out,
	output wire	gpio0_2_enable_vswitch_h,
	output wire	gpio0_2_enable_vdda_h,
	output wire	gpio0_2_vtrip_sel,
	output wire	gpio0_2_ib_mode_sel,
	output wire	gpio0_2_oe_n,
	input wire	gpio0_2_in_h,
	input wire	gpio0_2_zero,
	input wire	gpio0_2_one,
	input wire	gpio0_3_tie_lo_esd,
	input wire	gpio0_3_in,
	input wire	gpio0_3_tie_hi_esd,
	output wire	gpio0_3_enable_vddio,
	output wire	gpio0_3_slow,
	inout wire	gpio0_3_pad_a_esd_0_h,
	inout wire	gpio0_3_pad_a_esd_1_h,
	inout wire	gpio0_3_pad_a_noesd_h,
	output wire	gpio0_3_analog_en,
	output wire	gpio0_3_analog_pol,
	output wire	gpio0_3_inp_dis,
	output wire	gpio0_3_enable_inp_h,
	output wire	gpio0_3_enable_h,
	output wire	gpio0_3_hld_h_n,
	output wire	gpio0_3_analog_sel,
	output wire	[2:0]	gpio0_3_dm,
	output wire	gpio0_3_hld_ovr,
	output wire	gpio0_3_out,
	output wire	gpio0_3_enable_vswitch_h,
	output wire	gpio0_3_enable_vdda_h,
	output wire	gpio0_3_vtrip_sel,
	output wire	gpio0_3_ib_mode_sel,
	output wire	gpio0_3_oe_n,
	input wire	gpio0_3_in_h,
	input wire	gpio0_3_zero,
	input wire	gpio0_3_one,
	input wire	gpio0_4_tie_lo_esd,
	input wire	gpio0_4_in,
	input wire	gpio0_4_tie_hi_esd,
	output wire	gpio0_4_enable_vddio,
	output wire	gpio0_4_slow,
	inout wire	gpio0_4_pad_a_esd_0_h,
	inout wire	gpio0_4_pad_a_esd_1_h,
	inout wire	gpio0_4_pad_a_noesd_h,
	output wire	gpio0_4_analog_en,
	output wire	gpio0_4_analog_pol,
	output wire	gpio0_4_inp_dis,
	output wire	gpio0_4_enable_inp_h,
	output wire	gpio0_4_enable_h,
	output wire	gpio0_4_hld_h_n,
	output wire	gpio0_4_analog_sel,
	output wire	[2:0]	gpio0_4_dm,
	output wire	gpio0_4_hld_ovr,
	output wire	gpio0_4_out,
	output wire	gpio0_4_enable_vswitch_h,
	output wire	gpio0_4_enable_vdda_h,
	output wire	gpio0_4_vtrip_sel,
	output wire	gpio0_4_ib_mode_sel,
	output wire	gpio0_4_oe_n,
	input wire	gpio0_4_in_h,
	input wire	gpio0_4_zero,
	input wire	gpio0_4_one,
	input wire	gpio0_5_tie_lo_esd,
	input wire	gpio0_5_in,
	input wire	gpio0_5_tie_hi_esd,
	output wire	gpio0_5_enable_vddio,
	output wire	gpio0_5_slow,
	inout wire	gpio0_5_pad_a_esd_0_h,
	inout wire	gpio0_5_pad_a_esd_1_h,
	inout wire	gpio0_5_pad_a_noesd_h,
	output wire	gpio0_5_analog_en,
	output wire	gpio0_5_analog_pol,
	output wire	gpio0_5_inp_dis,
	output wire	gpio0_5_enable_inp_h,
	output wire	gpio0_5_enable_h,
	output wire	gpio0_5_hld_h_n,
	output wire	gpio0_5_analog_sel,
	output wire	[2:0]	gpio0_5_dm,
	output wire	gpio0_5_hld_ovr,
	output wire	gpio0_5_out,
	output wire	gpio0_5_enable_vswitch_h,
	output wire	gpio0_5_enable_vdda_h,
	output wire	gpio0_5_vtrip_sel,
	output wire	gpio0_5_ib_mode_sel,
	output wire	gpio0_5_oe_n,
	input wire	gpio0_5_in_h,
	input wire	gpio0_5_zero,
	input wire	gpio0_5_one,
	input wire	gpio0_6_tie_lo_esd,
	input wire	gpio0_6_in,
	input wire	gpio0_6_tie_hi_esd,
	output wire	gpio0_6_enable_vddio,
	output wire	gpio0_6_slow,
	inout wire	gpio0_6_pad_a_esd_0_h,
	inout wire	gpio0_6_pad_a_esd_1_h,
	inout wire	gpio0_6_pad_a_noesd_h,
	output wire	gpio0_6_analog_en,
	output wire	gpio0_6_analog_pol,
	output wire	gpio0_6_inp_dis,
	output wire	gpio0_6_enable_inp_h,
	output wire	gpio0_6_enable_h,
	output wire	gpio0_6_hld_h_n,
	output wire	gpio0_6_analog_sel,
	output wire	[2:0]	gpio0_6_dm,
	output wire	gpio0_6_hld_ovr,
	output wire	gpio0_6_out,
	output wire	gpio0_6_enable_vswitch_h,
	output wire	gpio0_6_enable_vdda_h,
	output wire	gpio0_6_vtrip_sel,
	output wire	gpio0_6_ib_mode_sel,
	output wire	gpio0_6_oe_n,
	input wire	gpio0_6_in_h,
	input wire	gpio0_6_zero,
	input wire	gpio0_6_one,
	input wire	gpio0_7_tie_lo_esd,
	input wire	gpio0_7_in,
	input wire	gpio0_7_tie_hi_esd,
	output wire	gpio0_7_enable_vddio,
	output wire	gpio0_7_slow,
	inout wire	gpio0_7_pad_a_esd_0_h,
	inout wire	gpio0_7_pad_a_esd_1_h,
	inout wire	gpio0_7_pad_a_noesd_h,
	output wire	gpio0_7_analog_en,
	output wire	gpio0_7_analog_pol,
	output wire	gpio0_7_inp_dis,
	output wire	gpio0_7_enable_inp_h,
	output wire	gpio0_7_enable_h,
	output wire	gpio0_7_hld_h_n,
	output wire	gpio0_7_analog_sel,
	output wire	[2:0]	gpio0_7_dm,
	output wire	gpio0_7_hld_ovr,
	output wire	gpio0_7_out,
	output wire	gpio0_7_enable_vswitch_h,
	output wire	gpio0_7_enable_vdda_h,
	output wire	gpio0_7_vtrip_sel,
	output wire	gpio0_7_ib_mode_sel,
	output wire	gpio0_7_oe_n,
	input wire	gpio0_7_in_h,
	input wire	gpio0_7_zero,
	input wire	gpio0_7_one,
	input wire	gpio1_0_tie_hi_esd,
	output wire	[2:0]	gpio1_0_dm,
	output wire	gpio1_0_slow,
	output wire	gpio1_0_oe_n,
	input wire	gpio1_0_tie_lo_esd,
	output wire	gpio1_0_inp_dis,
	output wire	gpio1_0_enable_vddio,
	output wire	gpio1_0_vtrip_sel,
	output wire	[1:0]	gpio1_0_ib_mode_sel,
	output wire	gpio1_0_out,
	output wire	[1:0]	gpio1_0_slew_ctl,
	output wire	gpio1_0_analog_pol,
	output wire	gpio1_0_analog_sel,
	output wire	gpio1_0_hys_trim,
	output wire	gpio1_0_hld_ovr,
	input wire	gpio1_0_in_h,
	output wire	gpio1_0_enable_h,
	input wire	gpio1_0_in,
	output wire	gpio1_0_hld_h_n,
	output wire	gpio1_0_enable_vdda_h,
	output wire	gpio1_0_analog_en,
	output wire	gpio1_0_enable_inp_h,
	output wire	gpio1_0_enable_vswitch_h,
	inout wire	gpio1_0_pad_a_noesd_h,
	inout wire	gpio1_0_pad_a_esd_0_h,
	inout wire	gpio1_0_pad_a_esd_1_h,
	input wire	gpio1_0_zero,
	input wire	gpio1_0_one,
	input wire	gpio1_1_tie_hi_esd,
	output wire	[2:0]	gpio1_1_dm,
	output wire	gpio1_1_slow,
	output wire	gpio1_1_oe_n,
	input wire	gpio1_1_tie_lo_esd,
	output wire	gpio1_1_inp_dis,
	output wire	gpio1_1_enable_vddio,
	output wire	gpio1_1_vtrip_sel,
	output wire	[1:0]	gpio1_1_ib_mode_sel,
	output wire	gpio1_1_out,
	output wire	[1:0]	gpio1_1_slew_ctl,
	output wire	gpio1_1_analog_pol,
	output wire	gpio1_1_analog_sel,
	output wire	gpio1_1_hys_trim,
	output wire	gpio1_1_hld_ovr,
	input wire	gpio1_1_in_h,
	output wire	gpio1_1_enable_h,
	input wire	gpio1_1_in,
	output wire	gpio1_1_hld_h_n,
	output wire	gpio1_1_enable_vdda_h,
	output wire	gpio1_1_analog_en,
	output wire	gpio1_1_enable_inp_h,
	output wire	gpio1_1_enable_vswitch_h,
	inout wire	gpio1_1_pad_a_noesd_h,
	inout wire	gpio1_1_pad_a_esd_0_h,
	inout wire	gpio1_1_pad_a_esd_1_h,
	input wire	gpio1_1_zero,
	input wire	gpio1_1_one,
	input wire	gpio1_2_tie_hi_esd,
	output wire	[2:0]	gpio1_2_dm,
	output wire	gpio1_2_slow,
	output wire	gpio1_2_oe_n,
	input wire	gpio1_2_tie_lo_esd,
	output wire	gpio1_2_inp_dis,
	output wire	gpio1_2_enable_vddio,
	output wire	gpio1_2_vtrip_sel,
	output wire	[1:0]	gpio1_2_ib_mode_sel,
	output wire	gpio1_2_out,
	output wire	[1:0]	gpio1_2_slew_ctl,
	output wire	gpio1_2_analog_pol,
	output wire	gpio1_2_analog_sel,
	output wire	gpio1_2_hys_trim,
	output wire	gpio1_2_hld_ovr,
	input wire	gpio1_2_in_h,
	output wire	gpio1_2_enable_h,
	input wire	gpio1_2_in,
	output wire	gpio1_2_hld_h_n,
	output wire	gpio1_2_enable_vdda_h,
	output wire	gpio1_2_analog_en,
	output wire	gpio1_2_enable_inp_h,
	output wire	gpio1_2_enable_vswitch_h,
	inout wire	gpio1_2_pad_a_noesd_h,
	inout wire	gpio1_2_pad_a_esd_0_h,
	inout wire	gpio1_2_pad_a_esd_1_h,
	input wire	gpio1_2_zero,
	input wire	gpio1_2_one,
	input wire	gpio1_3_tie_hi_esd,
	output wire	[2:0]	gpio1_3_dm,
	output wire	gpio1_3_slow,
	output wire	gpio1_3_oe_n,
	input wire	gpio1_3_tie_lo_esd,
	output wire	gpio1_3_inp_dis,
	output wire	gpio1_3_enable_vddio,
	output wire	gpio1_3_vtrip_sel,
	output wire	[1:0]	gpio1_3_ib_mode_sel,
	output wire	gpio1_3_out,
	output wire	[1:0]	gpio1_3_slew_ctl,
	output wire	gpio1_3_analog_pol,
	output wire	gpio1_3_analog_sel,
	output wire	gpio1_3_hys_trim,
	output wire	gpio1_3_hld_ovr,
	input wire	gpio1_3_in_h,
	output wire	gpio1_3_enable_h,
	input wire	gpio1_3_in,
	output wire	gpio1_3_hld_h_n,
	output wire	gpio1_3_enable_vdda_h,
	output wire	gpio1_3_analog_en,
	output wire	gpio1_3_enable_inp_h,
	output wire	gpio1_3_enable_vswitch_h,
	inout wire	gpio1_3_pad_a_noesd_h,
	inout wire	gpio1_3_pad_a_esd_0_h,
	inout wire	gpio1_3_pad_a_esd_1_h,
	input wire	gpio1_3_zero,
	input wire	gpio1_3_one,
	output wire	[4:0]	vref_e_ref_sel,
	inout wire	vref_e_vinref,
	output wire	vref_e_enable_h,
	output wire	vref_e_hld_h_n,
	output wire	vref_e_vrefgen_en,
	input wire	gpio1_4_tie_hi_esd,
	output wire	[2:0]	gpio1_4_dm,
	output wire	gpio1_4_slow,
	output wire	gpio1_4_oe_n,
	input wire	gpio1_4_tie_lo_esd,
	output wire	gpio1_4_inp_dis,
	output wire	gpio1_4_enable_vddio,
	output wire	gpio1_4_vtrip_sel,
	output wire	[1:0]	gpio1_4_ib_mode_sel,
	output wire	gpio1_4_out,
	output wire	[1:0]	gpio1_4_slew_ctl,
	output wire	gpio1_4_analog_pol,
	output wire	gpio1_4_analog_sel,
	output wire	gpio1_4_hys_trim,
	output wire	gpio1_4_hld_ovr,
	input wire	gpio1_4_in_h,
	output wire	gpio1_4_enable_h,
	input wire	gpio1_4_in,
	output wire	gpio1_4_hld_h_n,
	output wire	gpio1_4_enable_vdda_h,
	output wire	gpio1_4_analog_en,
	output wire	gpio1_4_enable_inp_h,
	output wire	gpio1_4_enable_vswitch_h,
	inout wire	gpio1_4_pad_a_noesd_h,
	inout wire	gpio1_4_pad_a_esd_0_h,
	inout wire	gpio1_4_pad_a_esd_1_h,
	input wire	gpio1_4_zero,
	input wire	gpio1_4_one,
	input wire	gpio1_5_tie_hi_esd,
	output wire	[2:0]	gpio1_5_dm,
	output wire	gpio1_5_slow,
	output wire	gpio1_5_oe_n,
	input wire	gpio1_5_tie_lo_esd,
	output wire	gpio1_5_inp_dis,
	output wire	gpio1_5_enable_vddio,
	output wire	gpio1_5_vtrip_sel,
	output wire	[1:0]	gpio1_5_ib_mode_sel,
	output wire	gpio1_5_out,
	output wire	[1:0]	gpio1_5_slew_ctl,
	output wire	gpio1_5_analog_pol,
	output wire	gpio1_5_analog_sel,
	output wire	gpio1_5_hys_trim,
	output wire	gpio1_5_hld_ovr,
	input wire	gpio1_5_in_h,
	output wire	gpio1_5_enable_h,
	input wire	gpio1_5_in,
	output wire	gpio1_5_hld_h_n,
	output wire	gpio1_5_enable_vdda_h,
	output wire	gpio1_5_analog_en,
	output wire	gpio1_5_enable_inp_h,
	output wire	gpio1_5_enable_vswitch_h,
	inout wire	gpio1_5_pad_a_noesd_h,
	inout wire	gpio1_5_pad_a_esd_0_h,
	inout wire	gpio1_5_pad_a_esd_1_h,
	input wire	gpio1_5_zero,
	input wire	gpio1_5_one,
	input wire	gpio1_6_tie_hi_esd,
	output wire	[2:0]	gpio1_6_dm,
	output wire	gpio1_6_slow,
	output wire	gpio1_6_oe_n,
	input wire	gpio1_6_tie_lo_esd,
	output wire	gpio1_6_inp_dis,
	output wire	gpio1_6_enable_vddio,
	output wire	gpio1_6_vtrip_sel,
	output wire	[1:0]	gpio1_6_ib_mode_sel,
	output wire	gpio1_6_out,
	output wire	[1:0]	gpio1_6_slew_ctl,
	output wire	gpio1_6_analog_pol,
	output wire	gpio1_6_analog_sel,
	output wire	gpio1_6_hys_trim,
	output wire	gpio1_6_hld_ovr,
	input wire	gpio1_6_in_h,
	output wire	gpio1_6_enable_h,
	input wire	gpio1_6_in,
	output wire	gpio1_6_hld_h_n,
	output wire	gpio1_6_enable_vdda_h,
	output wire	gpio1_6_analog_en,
	output wire	gpio1_6_enable_inp_h,
	output wire	gpio1_6_enable_vswitch_h,
	inout wire	gpio1_6_pad_a_noesd_h,
	inout wire	gpio1_6_pad_a_esd_0_h,
	inout wire	gpio1_6_pad_a_esd_1_h,
	input wire	gpio1_6_zero,
	input wire	gpio1_6_one,
	input wire	gpio1_7_tie_hi_esd,
	output wire	[2:0]	gpio1_7_dm,
	output wire	gpio1_7_slow,
	output wire	gpio1_7_oe_n,
	input wire	gpio1_7_tie_lo_esd,
	output wire	gpio1_7_inp_dis,
	output wire	gpio1_7_enable_vddio,
	output wire	gpio1_7_vtrip_sel,
	output wire	[1:0]	gpio1_7_ib_mode_sel,
	output wire	gpio1_7_out,
	output wire	[1:0]	gpio1_7_slew_ctl,
	output wire	gpio1_7_analog_pol,
	output wire	gpio1_7_analog_sel,
	output wire	gpio1_7_hys_trim,
	output wire	gpio1_7_hld_ovr,
	input wire	gpio1_7_in_h,
	output wire	gpio1_7_enable_h,
	input wire	gpio1_7_in,
	output wire	gpio1_7_hld_h_n,
	output wire	gpio1_7_enable_vdda_h,
	output wire	gpio1_7_analog_en,
	output wire	gpio1_7_enable_inp_h,
	output wire	gpio1_7_enable_vswitch_h,
	inout wire	gpio1_7_pad_a_noesd_h,
	inout wire	gpio1_7_pad_a_esd_0_h,
	inout wire	gpio1_7_pad_a_esd_1_h,
	input wire	gpio1_7_zero,
	input wire	gpio1_7_one,
	input wire	gpio2_0_tie_lo_esd,
	input wire	gpio2_0_in,
	input wire	gpio2_0_tie_hi_esd,
	output wire	gpio2_0_enable_vddio,
	output wire	gpio2_0_slow,
	inout wire	gpio2_0_pad_a_esd_0_h,
	inout wire	gpio2_0_pad_a_esd_1_h,
	inout wire	gpio2_0_pad_a_noesd_h,
	output wire	gpio2_0_analog_en,
	output wire	gpio2_0_analog_pol,
	output wire	gpio2_0_inp_dis,
	output wire	gpio2_0_enable_inp_h,
	output wire	gpio2_0_enable_h,
	output wire	gpio2_0_hld_h_n,
	output wire	gpio2_0_analog_sel,
	output wire	[2:0]	gpio2_0_dm,
	output wire	gpio2_0_hld_ovr,
	output wire	gpio2_0_out,
	output wire	gpio2_0_enable_vswitch_h,
	output wire	gpio2_0_enable_vdda_h,
	output wire	gpio2_0_vtrip_sel,
	output wire	gpio2_0_ib_mode_sel,
	output wire	gpio2_0_oe_n,
	input wire	gpio2_0_in_h,
	input wire	gpio2_0_zero,
	input wire	gpio2_0_one,
	input wire	gpio2_1_tie_lo_esd,
	input wire	gpio2_1_in,
	input wire	gpio2_1_tie_hi_esd,
	output wire	gpio2_1_enable_vddio,
	output wire	gpio2_1_slow,
	inout wire	gpio2_1_pad_a_esd_0_h,
	inout wire	gpio2_1_pad_a_esd_1_h,
	inout wire	gpio2_1_pad_a_noesd_h,
	output wire	gpio2_1_analog_en,
	output wire	gpio2_1_analog_pol,
	output wire	gpio2_1_inp_dis,
	output wire	gpio2_1_enable_inp_h,
	output wire	gpio2_1_enable_h,
	output wire	gpio2_1_hld_h_n,
	output wire	gpio2_1_analog_sel,
	output wire	[2:0]	gpio2_1_dm,
	output wire	gpio2_1_hld_ovr,
	output wire	gpio2_1_out,
	output wire	gpio2_1_enable_vswitch_h,
	output wire	gpio2_1_enable_vdda_h,
	output wire	gpio2_1_vtrip_sel,
	output wire	gpio2_1_ib_mode_sel,
	output wire	gpio2_1_oe_n,
	input wire	gpio2_1_in_h,
	input wire	gpio2_1_zero,
	input wire	gpio2_1_one,
	input wire	gpio2_2_tie_lo_esd,
	input wire	gpio2_2_in,
	input wire	gpio2_2_tie_hi_esd,
	output wire	gpio2_2_enable_vddio,
	output wire	gpio2_2_slow,
	inout wire	gpio2_2_pad_a_esd_0_h,
	inout wire	gpio2_2_pad_a_esd_1_h,
	inout wire	gpio2_2_pad_a_noesd_h,
	output wire	gpio2_2_analog_en,
	output wire	gpio2_2_analog_pol,
	output wire	gpio2_2_inp_dis,
	output wire	gpio2_2_enable_inp_h,
	output wire	gpio2_2_enable_h,
	output wire	gpio2_2_hld_h_n,
	output wire	gpio2_2_analog_sel,
	output wire	[2:0]	gpio2_2_dm,
	output wire	gpio2_2_hld_ovr,
	output wire	gpio2_2_out,
	output wire	gpio2_2_enable_vswitch_h,
	output wire	gpio2_2_enable_vdda_h,
	output wire	gpio2_2_vtrip_sel,
	output wire	gpio2_2_ib_mode_sel,
	output wire	gpio2_2_oe_n,
	input wire	gpio2_2_in_h,
	input wire	gpio2_2_zero,
	input wire	gpio2_2_one,
	input wire	gpio2_3_tie_lo_esd,
	input wire	gpio2_3_in,
	input wire	gpio2_3_tie_hi_esd,
	output wire	gpio2_3_enable_vddio,
	output wire	gpio2_3_slow,
	inout wire	gpio2_3_pad_a_esd_0_h,
	inout wire	gpio2_3_pad_a_esd_1_h,
	inout wire	gpio2_3_pad_a_noesd_h,
	output wire	gpio2_3_analog_en,
	output wire	gpio2_3_analog_pol,
	output wire	gpio2_3_inp_dis,
	output wire	gpio2_3_enable_inp_h,
	output wire	gpio2_3_enable_h,
	output wire	gpio2_3_hld_h_n,
	output wire	gpio2_3_analog_sel,
	output wire	[2:0]	gpio2_3_dm,
	output wire	gpio2_3_hld_ovr,
	output wire	gpio2_3_out,
	output wire	gpio2_3_enable_vswitch_h,
	output wire	gpio2_3_enable_vdda_h,
	output wire	gpio2_3_vtrip_sel,
	output wire	gpio2_3_ib_mode_sel,
	output wire	gpio2_3_oe_n,
	input wire	gpio2_3_in_h,
	input wire	gpio2_3_zero,
	input wire	gpio2_3_one,
	input wire	gpio2_4_tie_lo_esd,
	input wire	gpio2_4_in,
	input wire	gpio2_4_tie_hi_esd,
	output wire	gpio2_4_enable_vddio,
	output wire	gpio2_4_slow,
	inout wire	gpio2_4_pad_a_esd_0_h,
	inout wire	gpio2_4_pad_a_esd_1_h,
	inout wire	gpio2_4_pad_a_noesd_h,
	output wire	gpio2_4_analog_en,
	output wire	gpio2_4_analog_pol,
	output wire	gpio2_4_inp_dis,
	output wire	gpio2_4_enable_inp_h,
	output wire	gpio2_4_enable_h,
	output wire	gpio2_4_hld_h_n,
	output wire	gpio2_4_analog_sel,
	output wire	[2:0]	gpio2_4_dm,
	output wire	gpio2_4_hld_ovr,
	output wire	gpio2_4_out,
	output wire	gpio2_4_enable_vswitch_h,
	output wire	gpio2_4_enable_vdda_h,
	output wire	gpio2_4_vtrip_sel,
	output wire	gpio2_4_ib_mode_sel,
	output wire	gpio2_4_oe_n,
	input wire	gpio2_4_in_h,
	input wire	gpio2_4_zero,
	input wire	gpio2_4_one,
	input wire	gpio2_5_tie_lo_esd,
	input wire	gpio2_5_in,
	input wire	gpio2_5_tie_hi_esd,
	output wire	gpio2_5_enable_vddio,
	output wire	gpio2_5_slow,
	inout wire	gpio2_5_pad_a_esd_0_h,
	inout wire	gpio2_5_pad_a_esd_1_h,
	inout wire	gpio2_5_pad_a_noesd_h,
	output wire	gpio2_5_analog_en,
	output wire	gpio2_5_analog_pol,
	output wire	gpio2_5_inp_dis,
	output wire	gpio2_5_enable_inp_h,
	output wire	gpio2_5_enable_h,
	output wire	gpio2_5_hld_h_n,
	output wire	gpio2_5_analog_sel,
	output wire	[2:0]	gpio2_5_dm,
	output wire	gpio2_5_hld_ovr,
	output wire	gpio2_5_out,
	output wire	gpio2_5_enable_vswitch_h,
	output wire	gpio2_5_enable_vdda_h,
	output wire	gpio2_5_vtrip_sel,
	output wire	gpio2_5_ib_mode_sel,
	output wire	gpio2_5_oe_n,
	input wire	gpio2_5_in_h,
	input wire	gpio2_5_zero,
	input wire	gpio2_5_one,
	input wire	gpio2_6_tie_lo_esd,
	input wire	gpio2_6_in,
	input wire	gpio2_6_tie_hi_esd,
	output wire	gpio2_6_enable_vddio,
	output wire	gpio2_6_slow,
	inout wire	gpio2_6_pad_a_esd_0_h,
	inout wire	gpio2_6_pad_a_esd_1_h,
	inout wire	gpio2_6_pad_a_noesd_h,
	output wire	gpio2_6_analog_en,
	output wire	gpio2_6_analog_pol,
	output wire	gpio2_6_inp_dis,
	output wire	gpio2_6_enable_inp_h,
	output wire	gpio2_6_enable_h,
	output wire	gpio2_6_hld_h_n,
	output wire	gpio2_6_analog_sel,
	output wire	[2:0]	gpio2_6_dm,
	output wire	gpio2_6_hld_ovr,
	output wire	gpio2_6_out,
	output wire	gpio2_6_enable_vswitch_h,
	output wire	gpio2_6_enable_vdda_h,
	output wire	gpio2_6_vtrip_sel,
	output wire	gpio2_6_ib_mode_sel,
	output wire	gpio2_6_oe_n,
	input wire	gpio2_6_in_h,
	input wire	gpio2_6_zero,
	input wire	gpio2_6_one,
	input wire	gpio2_7_tie_lo_esd,
	input wire	gpio2_7_in,
	input wire	gpio2_7_tie_hi_esd,
	output wire	gpio2_7_enable_vddio,
	output wire	gpio2_7_slow,
	inout wire	gpio2_7_pad_a_esd_0_h,
	inout wire	gpio2_7_pad_a_esd_1_h,
	inout wire	gpio2_7_pad_a_noesd_h,
	output wire	gpio2_7_analog_en,
	output wire	gpio2_7_analog_pol,
	output wire	gpio2_7_inp_dis,
	output wire	gpio2_7_enable_inp_h,
	output wire	gpio2_7_enable_h,
	output wire	gpio2_7_hld_h_n,
	output wire	gpio2_7_analog_sel,
	output wire	[2:0]	gpio2_7_dm,
	output wire	gpio2_7_hld_ovr,
	output wire	gpio2_7_out,
	output wire	gpio2_7_enable_vswitch_h,
	output wire	gpio2_7_enable_vdda_h,
	output wire	gpio2_7_vtrip_sel,
	output wire	gpio2_7_ib_mode_sel,
	output wire	gpio2_7_oe_n,
	input wire	gpio2_7_in_h,
	input wire	gpio2_7_zero,
	input wire	gpio2_7_one,
	output wire	muxsplit_ne_hld_vdda_h_n,
	output wire	muxsplit_ne_enable_vdda_h,
	output wire	muxsplit_ne_switch_aa_sl,
	output wire	muxsplit_ne_switch_aa_s0,
	output wire	muxsplit_ne_switch_bb_s0,
	output wire	muxsplit_ne_switch_bb_sl,
	output wire	muxsplit_ne_switch_bb_sr,
	output wire	muxsplit_ne_switch_aa_sr,
	input wire	gpio3_0_tie_lo_esd,
	input wire	gpio3_0_in,
	input wire	gpio3_0_tie_hi_esd,
	output wire	gpio3_0_enable_vddio,
	output wire	gpio3_0_slow,
	inout wire	gpio3_0_pad_a_esd_0_h,
	inout wire	gpio3_0_pad_a_esd_1_h,
	inout wire	gpio3_0_pad_a_noesd_h,
	output wire	gpio3_0_analog_en,
	output wire	gpio3_0_analog_pol,
	output wire	gpio3_0_inp_dis,
	output wire	gpio3_0_enable_inp_h,
	output wire	gpio3_0_enable_h,
	output wire	gpio3_0_hld_h_n,
	output wire	gpio3_0_analog_sel,
	output wire	[2:0]	gpio3_0_dm,
	output wire	gpio3_0_hld_ovr,
	output wire	gpio3_0_out,
	output wire	gpio3_0_enable_vswitch_h,
	output wire	gpio3_0_enable_vdda_h,
	output wire	gpio3_0_vtrip_sel,
	output wire	gpio3_0_ib_mode_sel,
	output wire	gpio3_0_oe_n,
	input wire	gpio3_0_in_h,
	input wire	gpio3_0_zero,
	input wire	gpio3_0_one,
	input wire	gpio3_1_tie_lo_esd,
	input wire	gpio3_1_in,
	input wire	gpio3_1_tie_hi_esd,
	output wire	gpio3_1_enable_vddio,
	output wire	gpio3_1_slow,
	inout wire	gpio3_1_pad_a_esd_0_h,
	inout wire	gpio3_1_pad_a_esd_1_h,
	inout wire	gpio3_1_pad_a_noesd_h,
	output wire	gpio3_1_analog_en,
	output wire	gpio3_1_analog_pol,
	output wire	gpio3_1_inp_dis,
	output wire	gpio3_1_enable_inp_h,
	output wire	gpio3_1_enable_h,
	output wire	gpio3_1_hld_h_n,
	output wire	gpio3_1_analog_sel,
	output wire	[2:0]	gpio3_1_dm,
	output wire	gpio3_1_hld_ovr,
	output wire	gpio3_1_out,
	output wire	gpio3_1_enable_vswitch_h,
	output wire	gpio3_1_enable_vdda_h,
	output wire	gpio3_1_vtrip_sel,
	output wire	gpio3_1_ib_mode_sel,
	output wire	gpio3_1_oe_n,
	input wire	gpio3_1_in_h,
	input wire	gpio3_1_zero,
	input wire	gpio3_1_one,
	input wire	gpio3_2_tie_lo_esd,
	input wire	gpio3_2_in,
	input wire	gpio3_2_tie_hi_esd,
	output wire	gpio3_2_enable_vddio,
	output wire	gpio3_2_slow,
	inout wire	gpio3_2_pad_a_esd_0_h,
	inout wire	gpio3_2_pad_a_esd_1_h,
	inout wire	gpio3_2_pad_a_noesd_h,
	output wire	gpio3_2_analog_en,
	output wire	gpio3_2_analog_pol,
	output wire	gpio3_2_inp_dis,
	output wire	gpio3_2_enable_inp_h,
	output wire	gpio3_2_enable_h,
	output wire	gpio3_2_hld_h_n,
	output wire	gpio3_2_analog_sel,
	output wire	[2:0]	gpio3_2_dm,
	output wire	gpio3_2_hld_ovr,
	output wire	gpio3_2_out,
	output wire	gpio3_2_enable_vswitch_h,
	output wire	gpio3_2_enable_vdda_h,
	output wire	gpio3_2_vtrip_sel,
	output wire	gpio3_2_ib_mode_sel,
	output wire	gpio3_2_oe_n,
	input wire	gpio3_2_in_h,
	input wire	gpio3_2_zero,
	input wire	gpio3_2_one,
	input wire	gpio3_3_tie_lo_esd,
	input wire	gpio3_3_in,
	input wire	gpio3_3_tie_hi_esd,
	output wire	gpio3_3_enable_vddio,
	output wire	gpio3_3_slow,
	inout wire	gpio3_3_pad_a_esd_0_h,
	inout wire	gpio3_3_pad_a_esd_1_h,
	inout wire	gpio3_3_pad_a_noesd_h,
	output wire	gpio3_3_analog_en,
	output wire	gpio3_3_analog_pol,
	output wire	gpio3_3_inp_dis,
	output wire	gpio3_3_enable_inp_h,
	output wire	gpio3_3_enable_h,
	output wire	gpio3_3_hld_h_n,
	output wire	gpio3_3_analog_sel,
	output wire	[2:0]	gpio3_3_dm,
	output wire	gpio3_3_hld_ovr,
	output wire	gpio3_3_out,
	output wire	gpio3_3_enable_vswitch_h,
	output wire	gpio3_3_enable_vdda_h,
	output wire	gpio3_3_vtrip_sel,
	output wire	gpio3_3_ib_mode_sel,
	output wire	gpio3_3_oe_n,
	input wire	gpio3_3_in_h,
	input wire	gpio3_3_zero,
	input wire	gpio3_3_one,
	input wire	gpio3_4_tie_lo_esd,
	input wire	gpio3_4_in,
	input wire	gpio3_4_tie_hi_esd,
	output wire	gpio3_4_enable_vddio,
	output wire	gpio3_4_slow,
	inout wire	gpio3_4_pad_a_esd_0_h,
	inout wire	gpio3_4_pad_a_esd_1_h,
	inout wire	gpio3_4_pad_a_noesd_h,
	output wire	gpio3_4_analog_en,
	output wire	gpio3_4_analog_pol,
	output wire	gpio3_4_inp_dis,
	output wire	gpio3_4_enable_inp_h,
	output wire	gpio3_4_enable_h,
	output wire	gpio3_4_hld_h_n,
	output wire	gpio3_4_analog_sel,
	output wire	[2:0]	gpio3_4_dm,
	output wire	gpio3_4_hld_ovr,
	output wire	gpio3_4_out,
	output wire	gpio3_4_enable_vswitch_h,
	output wire	gpio3_4_enable_vdda_h,
	output wire	gpio3_4_vtrip_sel,
	output wire	gpio3_4_ib_mode_sel,
	output wire	gpio3_4_oe_n,
	input wire	gpio3_4_in_h,
	input wire	gpio3_4_zero,
	input wire	gpio3_4_one,
	input wire	gpio3_5_tie_lo_esd,
	input wire	gpio3_5_in,
	input wire	gpio3_5_tie_hi_esd,
	output wire	gpio3_5_enable_vddio,
	output wire	gpio3_5_slow,
	inout wire	gpio3_5_pad_a_esd_0_h,
	inout wire	gpio3_5_pad_a_esd_1_h,
	inout wire	gpio3_5_pad_a_noesd_h,
	output wire	gpio3_5_analog_en,
	output wire	gpio3_5_analog_pol,
	output wire	gpio3_5_inp_dis,
	output wire	gpio3_5_enable_inp_h,
	output wire	gpio3_5_enable_h,
	output wire	gpio3_5_hld_h_n,
	output wire	gpio3_5_analog_sel,
	output wire	[2:0]	gpio3_5_dm,
	output wire	gpio3_5_hld_ovr,
	output wire	gpio3_5_out,
	output wire	gpio3_5_enable_vswitch_h,
	output wire	gpio3_5_enable_vdda_h,
	output wire	gpio3_5_vtrip_sel,
	output wire	gpio3_5_ib_mode_sel,
	output wire	gpio3_5_oe_n,
	input wire	gpio3_5_in_h,
	input wire	gpio3_5_zero,
	input wire	gpio3_5_one,
	input wire	gpio3_6_tie_lo_esd,
	input wire	gpio3_6_in,
	input wire	gpio3_6_tie_hi_esd,
	output wire	gpio3_6_enable_vddio,
	output wire	gpio3_6_slow,
	inout wire	gpio3_6_pad_a_esd_0_h,
	inout wire	gpio3_6_pad_a_esd_1_h,
	inout wire	gpio3_6_pad_a_noesd_h,
	output wire	gpio3_6_analog_en,
	output wire	gpio3_6_analog_pol,
	output wire	gpio3_6_inp_dis,
	output wire	gpio3_6_enable_inp_h,
	output wire	gpio3_6_enable_h,
	output wire	gpio3_6_hld_h_n,
	output wire	gpio3_6_analog_sel,
	output wire	[2:0]	gpio3_6_dm,
	output wire	gpio3_6_hld_ovr,
	output wire	gpio3_6_out,
	output wire	gpio3_6_enable_vswitch_h,
	output wire	gpio3_6_enable_vdda_h,
	output wire	gpio3_6_vtrip_sel,
	output wire	gpio3_6_ib_mode_sel,
	output wire	gpio3_6_oe_n,
	input wire	gpio3_6_in_h,
	input wire	gpio3_6_zero,
	input wire	gpio3_6_one,
	input wire	gpio3_7_tie_lo_esd,
	input wire	gpio3_7_in,
	input wire	gpio3_7_tie_hi_esd,
	output wire	gpio3_7_enable_vddio,
	output wire	gpio3_7_slow,
	inout wire	gpio3_7_pad_a_esd_0_h,
	inout wire	gpio3_7_pad_a_esd_1_h,
	inout wire	gpio3_7_pad_a_noesd_h,
	output wire	gpio3_7_analog_en,
	output wire	gpio3_7_analog_pol,
	output wire	gpio3_7_inp_dis,
	output wire	gpio3_7_enable_inp_h,
	output wire	gpio3_7_enable_h,
	output wire	gpio3_7_hld_h_n,
	output wire	gpio3_7_analog_sel,
	output wire	[2:0]	gpio3_7_dm,
	output wire	gpio3_7_hld_ovr,
	output wire	gpio3_7_out,
	output wire	gpio3_7_enable_vswitch_h,
	output wire	gpio3_7_enable_vdda_h,
	output wire	gpio3_7_vtrip_sel,
	output wire	gpio3_7_ib_mode_sel,
	output wire	gpio3_7_oe_n,
	input wire	gpio3_7_in_h,
	input wire	gpio3_7_zero,
	input wire	gpio3_7_one,
	inout wire	analog_0_core,
	inout wire	analog_1_core,
	input wire	gpio4_0_tie_lo_esd,
	input wire	gpio4_0_in,
	input wire	gpio4_0_tie_hi_esd,
	output wire	gpio4_0_enable_vddio,
	output wire	gpio4_0_slow,
	inout wire	gpio4_0_pad_a_esd_0_h,
	inout wire	gpio4_0_pad_a_esd_1_h,
	inout wire	gpio4_0_pad_a_noesd_h,
	output wire	gpio4_0_analog_en,
	output wire	gpio4_0_analog_pol,
	output wire	gpio4_0_inp_dis,
	output wire	gpio4_0_enable_inp_h,
	output wire	gpio4_0_enable_h,
	output wire	gpio4_0_hld_h_n,
	output wire	gpio4_0_analog_sel,
	output wire	[2:0]	gpio4_0_dm,
	output wire	gpio4_0_hld_ovr,
	output wire	gpio4_0_out,
	output wire	gpio4_0_enable_vswitch_h,
	output wire	gpio4_0_enable_vdda_h,
	output wire	gpio4_0_vtrip_sel,
	output wire	gpio4_0_ib_mode_sel,
	output wire	gpio4_0_oe_n,
	input wire	gpio4_0_in_h,
	input wire	gpio4_0_zero,
	input wire	gpio4_0_one,
	input wire	gpio4_1_tie_lo_esd,
	input wire	gpio4_1_in,
	input wire	gpio4_1_tie_hi_esd,
	output wire	gpio4_1_enable_vddio,
	output wire	gpio4_1_slow,
	inout wire	gpio4_1_pad_a_esd_0_h,
	inout wire	gpio4_1_pad_a_esd_1_h,
	inout wire	gpio4_1_pad_a_noesd_h,
	output wire	gpio4_1_analog_en,
	output wire	gpio4_1_analog_pol,
	output wire	gpio4_1_inp_dis,
	output wire	gpio4_1_enable_inp_h,
	output wire	gpio4_1_enable_h,
	output wire	gpio4_1_hld_h_n,
	output wire	gpio4_1_analog_sel,
	output wire	[2:0]	gpio4_1_dm,
	output wire	gpio4_1_hld_ovr,
	output wire	gpio4_1_out,
	output wire	gpio4_1_enable_vswitch_h,
	output wire	gpio4_1_enable_vdda_h,
	output wire	gpio4_1_vtrip_sel,
	output wire	gpio4_1_ib_mode_sel,
	output wire	gpio4_1_oe_n,
	input wire	gpio4_1_in_h,
	input wire	gpio4_1_zero,
	input wire	gpio4_1_one,
	input wire	gpio4_2_tie_lo_esd,
	input wire	gpio4_2_in,
	input wire	gpio4_2_tie_hi_esd,
	output wire	gpio4_2_enable_vddio,
	output wire	gpio4_2_slow,
	inout wire	gpio4_2_pad_a_esd_0_h,
	inout wire	gpio4_2_pad_a_esd_1_h,
	inout wire	gpio4_2_pad_a_noesd_h,
	output wire	gpio4_2_analog_en,
	output wire	gpio4_2_analog_pol,
	output wire	gpio4_2_inp_dis,
	output wire	gpio4_2_enable_inp_h,
	output wire	gpio4_2_enable_h,
	output wire	gpio4_2_hld_h_n,
	output wire	gpio4_2_analog_sel,
	output wire	[2:0]	gpio4_2_dm,
	output wire	gpio4_2_hld_ovr,
	output wire	gpio4_2_out,
	output wire	gpio4_2_enable_vswitch_h,
	output wire	gpio4_2_enable_vdda_h,
	output wire	gpio4_2_vtrip_sel,
	output wire	gpio4_2_ib_mode_sel,
	output wire	gpio4_2_oe_n,
	input wire	gpio4_2_in_h,
	input wire	gpio4_2_zero,
	input wire	gpio4_2_one,
	input wire	gpio4_3_tie_lo_esd,
	input wire	gpio4_3_in,
	input wire	gpio4_3_tie_hi_esd,
	output wire	gpio4_3_enable_vddio,
	output wire	gpio4_3_slow,
	inout wire	gpio4_3_pad_a_esd_0_h,
	inout wire	gpio4_3_pad_a_esd_1_h,
	inout wire	gpio4_3_pad_a_noesd_h,
	output wire	gpio4_3_analog_en,
	output wire	gpio4_3_analog_pol,
	output wire	gpio4_3_inp_dis,
	output wire	gpio4_3_enable_inp_h,
	output wire	gpio4_3_enable_h,
	output wire	gpio4_3_hld_h_n,
	output wire	gpio4_3_analog_sel,
	output wire	[2:0]	gpio4_3_dm,
	output wire	gpio4_3_hld_ovr,
	output wire	gpio4_3_out,
	output wire	gpio4_3_enable_vswitch_h,
	output wire	gpio4_3_enable_vdda_h,
	output wire	gpio4_3_vtrip_sel,
	output wire	gpio4_3_ib_mode_sel,
	output wire	gpio4_3_oe_n,
	input wire	gpio4_3_in_h,
	input wire	gpio4_3_zero,
	input wire	gpio4_3_one,
	input wire	gpio4_4_tie_lo_esd,
	input wire	gpio4_4_in,
	input wire	gpio4_4_tie_hi_esd,
	output wire	gpio4_4_enable_vddio,
	output wire	gpio4_4_slow,
	inout wire	gpio4_4_pad_a_esd_0_h,
	inout wire	gpio4_4_pad_a_esd_1_h,
	inout wire	gpio4_4_pad_a_noesd_h,
	output wire	gpio4_4_analog_en,
	output wire	gpio4_4_analog_pol,
	output wire	gpio4_4_inp_dis,
	output wire	gpio4_4_enable_inp_h,
	output wire	gpio4_4_enable_h,
	output wire	gpio4_4_hld_h_n,
	output wire	gpio4_4_analog_sel,
	output wire	[2:0]	gpio4_4_dm,
	output wire	gpio4_4_hld_ovr,
	output wire	gpio4_4_out,
	output wire	gpio4_4_enable_vswitch_h,
	output wire	gpio4_4_enable_vdda_h,
	output wire	gpio4_4_vtrip_sel,
	output wire	gpio4_4_ib_mode_sel,
	output wire	gpio4_4_oe_n,
	input wire	gpio4_4_in_h,
	input wire	gpio4_4_zero,
	input wire	gpio4_4_one,
	input wire	gpio4_5_tie_lo_esd,
	input wire	gpio4_5_in,
	input wire	gpio4_5_tie_hi_esd,
	output wire	gpio4_5_enable_vddio,
	output wire	gpio4_5_slow,
	inout wire	gpio4_5_pad_a_esd_0_h,
	inout wire	gpio4_5_pad_a_esd_1_h,
	inout wire	gpio4_5_pad_a_noesd_h,
	output wire	gpio4_5_analog_en,
	output wire	gpio4_5_analog_pol,
	output wire	gpio4_5_inp_dis,
	output wire	gpio4_5_enable_inp_h,
	output wire	gpio4_5_enable_h,
	output wire	gpio4_5_hld_h_n,
	output wire	gpio4_5_analog_sel,
	output wire	[2:0]	gpio4_5_dm,
	output wire	gpio4_5_hld_ovr,
	output wire	gpio4_5_out,
	output wire	gpio4_5_enable_vswitch_h,
	output wire	gpio4_5_enable_vdda_h,
	output wire	gpio4_5_vtrip_sel,
	output wire	gpio4_5_ib_mode_sel,
	output wire	gpio4_5_oe_n,
	input wire	gpio4_5_in_h,
	input wire	gpio4_5_zero,
	input wire	gpio4_5_one,
	input wire	gpio4_6_tie_lo_esd,
	input wire	gpio4_6_in,
	input wire	gpio4_6_tie_hi_esd,
	output wire	gpio4_6_enable_vddio,
	output wire	gpio4_6_slow,
	inout wire	gpio4_6_pad_a_esd_0_h,
	inout wire	gpio4_6_pad_a_esd_1_h,
	inout wire	gpio4_6_pad_a_noesd_h,
	output wire	gpio4_6_analog_en,
	output wire	gpio4_6_analog_pol,
	output wire	gpio4_6_inp_dis,
	output wire	gpio4_6_enable_inp_h,
	output wire	gpio4_6_enable_h,
	output wire	gpio4_6_hld_h_n,
	output wire	gpio4_6_analog_sel,
	output wire	[2:0]	gpio4_6_dm,
	output wire	gpio4_6_hld_ovr,
	output wire	gpio4_6_out,
	output wire	gpio4_6_enable_vswitch_h,
	output wire	gpio4_6_enable_vdda_h,
	output wire	gpio4_6_vtrip_sel,
	output wire	gpio4_6_ib_mode_sel,
	output wire	gpio4_6_oe_n,
	input wire	gpio4_6_in_h,
	input wire	gpio4_6_zero,
	input wire	gpio4_6_one,
	input wire	gpio4_7_tie_lo_esd,
	input wire	gpio4_7_in,
	input wire	gpio4_7_tie_hi_esd,
	output wire	gpio4_7_enable_vddio,
	output wire	gpio4_7_slow,
	inout wire	gpio4_7_pad_a_esd_0_h,
	inout wire	gpio4_7_pad_a_esd_1_h,
	inout wire	gpio4_7_pad_a_noesd_h,
	output wire	gpio4_7_analog_en,
	output wire	gpio4_7_analog_pol,
	output wire	gpio4_7_inp_dis,
	output wire	gpio4_7_enable_inp_h,
	output wire	gpio4_7_enable_h,
	output wire	gpio4_7_hld_h_n,
	output wire	gpio4_7_analog_sel,
	output wire	[2:0]	gpio4_7_dm,
	output wire	gpio4_7_hld_ovr,
	output wire	gpio4_7_out,
	output wire	gpio4_7_enable_vswitch_h,
	output wire	gpio4_7_enable_vdda_h,
	output wire	gpio4_7_vtrip_sel,
	output wire	gpio4_7_ib_mode_sel,
	output wire	gpio4_7_oe_n,
	input wire	gpio4_7_in_h,
	input wire	gpio4_7_zero,
	input wire	gpio4_7_one,
	output wire	muxsplit_nw_hld_vdda_h_n,
	output wire	muxsplit_nw_enable_vdda_h,
	output wire	muxsplit_nw_switch_aa_sl,
	output wire	muxsplit_nw_switch_aa_s0,
	output wire	muxsplit_nw_switch_bb_s0,
	output wire	muxsplit_nw_switch_bb_sl,
	output wire	muxsplit_nw_switch_bb_sr,
	output wire	muxsplit_nw_switch_aa_sr,
	input wire	gpio5_0_tie_lo_esd,
	input wire	gpio5_0_in,
	input wire	gpio5_0_tie_hi_esd,
	output wire	gpio5_0_enable_vddio,
	output wire	gpio5_0_slow,
	inout wire	gpio5_0_pad_a_esd_0_h,
	inout wire	gpio5_0_pad_a_esd_1_h,
	inout wire	gpio5_0_pad_a_noesd_h,
	output wire	gpio5_0_analog_en,
	output wire	gpio5_0_analog_pol,
	output wire	gpio5_0_inp_dis,
	output wire	gpio5_0_enable_inp_h,
	output wire	gpio5_0_enable_h,
	output wire	gpio5_0_hld_h_n,
	output wire	gpio5_0_analog_sel,
	output wire	[2:0]	gpio5_0_dm,
	output wire	gpio5_0_hld_ovr,
	output wire	gpio5_0_out,
	output wire	gpio5_0_enable_vswitch_h,
	output wire	gpio5_0_enable_vdda_h,
	output wire	gpio5_0_vtrip_sel,
	output wire	gpio5_0_ib_mode_sel,
	output wire	gpio5_0_oe_n,
	input wire	gpio5_0_in_h,
	input wire	gpio5_0_zero,
	input wire	gpio5_0_one,
	input wire	gpio5_1_tie_lo_esd,
	input wire	gpio5_1_in,
	input wire	gpio5_1_tie_hi_esd,
	output wire	gpio5_1_enable_vddio,
	output wire	gpio5_1_slow,
	inout wire	gpio5_1_pad_a_esd_0_h,
	inout wire	gpio5_1_pad_a_esd_1_h,
	inout wire	gpio5_1_pad_a_noesd_h,
	output wire	gpio5_1_analog_en,
	output wire	gpio5_1_analog_pol,
	output wire	gpio5_1_inp_dis,
	output wire	gpio5_1_enable_inp_h,
	output wire	gpio5_1_enable_h,
	output wire	gpio5_1_hld_h_n,
	output wire	gpio5_1_analog_sel,
	output wire	[2:0]	gpio5_1_dm,
	output wire	gpio5_1_hld_ovr,
	output wire	gpio5_1_out,
	output wire	gpio5_1_enable_vswitch_h,
	output wire	gpio5_1_enable_vdda_h,
	output wire	gpio5_1_vtrip_sel,
	output wire	gpio5_1_ib_mode_sel,
	output wire	gpio5_1_oe_n,
	input wire	gpio5_1_in_h,
	input wire	gpio5_1_zero,
	input wire	gpio5_1_one,
	input wire	gpio5_2_tie_lo_esd,
	input wire	gpio5_2_in,
	input wire	gpio5_2_tie_hi_esd,
	output wire	gpio5_2_enable_vddio,
	output wire	gpio5_2_slow,
	inout wire	gpio5_2_pad_a_esd_0_h,
	inout wire	gpio5_2_pad_a_esd_1_h,
	inout wire	gpio5_2_pad_a_noesd_h,
	output wire	gpio5_2_analog_en,
	output wire	gpio5_2_analog_pol,
	output wire	gpio5_2_inp_dis,
	output wire	gpio5_2_enable_inp_h,
	output wire	gpio5_2_enable_h,
	output wire	gpio5_2_hld_h_n,
	output wire	gpio5_2_analog_sel,
	output wire	[2:0]	gpio5_2_dm,
	output wire	gpio5_2_hld_ovr,
	output wire	gpio5_2_out,
	output wire	gpio5_2_enable_vswitch_h,
	output wire	gpio5_2_enable_vdda_h,
	output wire	gpio5_2_vtrip_sel,
	output wire	gpio5_2_ib_mode_sel,
	output wire	gpio5_2_oe_n,
	input wire	gpio5_2_in_h,
	input wire	gpio5_2_zero,
	input wire	gpio5_2_one,
	input wire	gpio5_3_tie_lo_esd,
	input wire	gpio5_3_in,
	input wire	gpio5_3_tie_hi_esd,
	output wire	gpio5_3_enable_vddio,
	output wire	gpio5_3_slow,
	inout wire	gpio5_3_pad_a_esd_0_h,
	inout wire	gpio5_3_pad_a_esd_1_h,
	inout wire	gpio5_3_pad_a_noesd_h,
	output wire	gpio5_3_analog_en,
	output wire	gpio5_3_analog_pol,
	output wire	gpio5_3_inp_dis,
	output wire	gpio5_3_enable_inp_h,
	output wire	gpio5_3_enable_h,
	output wire	gpio5_3_hld_h_n,
	output wire	gpio5_3_analog_sel,
	output wire	[2:0]	gpio5_3_dm,
	output wire	gpio5_3_hld_ovr,
	output wire	gpio5_3_out,
	output wire	gpio5_3_enable_vswitch_h,
	output wire	gpio5_3_enable_vdda_h,
	output wire	gpio5_3_vtrip_sel,
	output wire	gpio5_3_ib_mode_sel,
	output wire	gpio5_3_oe_n,
	input wire	gpio5_3_in_h,
	input wire	gpio5_3_zero,
	input wire	gpio5_3_one,
	input wire	gpio5_4_tie_lo_esd,
	input wire	gpio5_4_in,
	input wire	gpio5_4_tie_hi_esd,
	output wire	gpio5_4_enable_vddio,
	output wire	gpio5_4_slow,
	inout wire	gpio5_4_pad_a_esd_0_h,
	inout wire	gpio5_4_pad_a_esd_1_h,
	inout wire	gpio5_4_pad_a_noesd_h,
	output wire	gpio5_4_analog_en,
	output wire	gpio5_4_analog_pol,
	output wire	gpio5_4_inp_dis,
	output wire	gpio5_4_enable_inp_h,
	output wire	gpio5_4_enable_h,
	output wire	gpio5_4_hld_h_n,
	output wire	gpio5_4_analog_sel,
	output wire	[2:0]	gpio5_4_dm,
	output wire	gpio5_4_hld_ovr,
	output wire	gpio5_4_out,
	output wire	gpio5_4_enable_vswitch_h,
	output wire	gpio5_4_enable_vdda_h,
	output wire	gpio5_4_vtrip_sel,
	output wire	gpio5_4_ib_mode_sel,
	output wire	gpio5_4_oe_n,
	input wire	gpio5_4_in_h,
	input wire	gpio5_4_zero,
	input wire	gpio5_4_one,
	input wire	gpio5_5_tie_lo_esd,
	input wire	gpio5_5_in,
	input wire	gpio5_5_tie_hi_esd,
	output wire	gpio5_5_enable_vddio,
	output wire	gpio5_5_slow,
	inout wire	gpio5_5_pad_a_esd_0_h,
	inout wire	gpio5_5_pad_a_esd_1_h,
	inout wire	gpio5_5_pad_a_noesd_h,
	output wire	gpio5_5_analog_en,
	output wire	gpio5_5_analog_pol,
	output wire	gpio5_5_inp_dis,
	output wire	gpio5_5_enable_inp_h,
	output wire	gpio5_5_enable_h,
	output wire	gpio5_5_hld_h_n,
	output wire	gpio5_5_analog_sel,
	output wire	[2:0]	gpio5_5_dm,
	output wire	gpio5_5_hld_ovr,
	output wire	gpio5_5_out,
	output wire	gpio5_5_enable_vswitch_h,
	output wire	gpio5_5_enable_vdda_h,
	output wire	gpio5_5_vtrip_sel,
	output wire	gpio5_5_ib_mode_sel,
	output wire	gpio5_5_oe_n,
	input wire	gpio5_5_in_h,
	input wire	gpio5_5_zero,
	input wire	gpio5_5_one,
	input wire	gpio5_6_tie_lo_esd,
	input wire	gpio5_6_in,
	input wire	gpio5_6_tie_hi_esd,
	output wire	gpio5_6_enable_vddio,
	output wire	gpio5_6_slow,
	inout wire	gpio5_6_pad_a_esd_0_h,
	inout wire	gpio5_6_pad_a_esd_1_h,
	inout wire	gpio5_6_pad_a_noesd_h,
	output wire	gpio5_6_analog_en,
	output wire	gpio5_6_analog_pol,
	output wire	gpio5_6_inp_dis,
	output wire	gpio5_6_enable_inp_h,
	output wire	gpio5_6_enable_h,
	output wire	gpio5_6_hld_h_n,
	output wire	gpio5_6_analog_sel,
	output wire	[2:0]	gpio5_6_dm,
	output wire	gpio5_6_hld_ovr,
	output wire	gpio5_6_out,
	output wire	gpio5_6_enable_vswitch_h,
	output wire	gpio5_6_enable_vdda_h,
	output wire	gpio5_6_vtrip_sel,
	output wire	gpio5_6_ib_mode_sel,
	output wire	gpio5_6_oe_n,
	input wire	gpio5_6_in_h,
	input wire	gpio5_6_zero,
	input wire	gpio5_6_one,
	input wire	gpio5_7_tie_lo_esd,
	input wire	gpio5_7_in,
	input wire	gpio5_7_tie_hi_esd,
	output wire	gpio5_7_enable_vddio,
	output wire	gpio5_7_slow,
	inout wire	gpio5_7_pad_a_esd_0_h,
	inout wire	gpio5_7_pad_a_esd_1_h,
	inout wire	gpio5_7_pad_a_noesd_h,
	output wire	gpio5_7_analog_en,
	output wire	gpio5_7_analog_pol,
	output wire	gpio5_7_inp_dis,
	output wire	gpio5_7_enable_inp_h,
	output wire	gpio5_7_enable_h,
	output wire	gpio5_7_hld_h_n,
	output wire	gpio5_7_analog_sel,
	output wire	[2:0]	gpio5_7_dm,
	output wire	gpio5_7_hld_ovr,
	output wire	gpio5_7_out,
	output wire	gpio5_7_enable_vswitch_h,
	output wire	gpio5_7_enable_vdda_h,
	output wire	gpio5_7_vtrip_sel,
	output wire	gpio5_7_ib_mode_sel,
	output wire	gpio5_7_oe_n,
	input wire	gpio5_7_in_h,
	input wire	gpio5_7_zero,
	input wire	gpio5_7_one,
	input wire	gpio6_0_tie_hi_esd,
	output wire	[2:0]	gpio6_0_dm,
	output wire	gpio6_0_slow,
	output wire	gpio6_0_oe_n,
	input wire	gpio6_0_tie_lo_esd,
	output wire	gpio6_0_inp_dis,
	output wire	gpio6_0_enable_vddio,
	output wire	gpio6_0_vtrip_sel,
	output wire	[1:0]	gpio6_0_ib_mode_sel,
	output wire	gpio6_0_out,
	output wire	[1:0]	gpio6_0_slew_ctl,
	output wire	gpio6_0_analog_pol,
	output wire	gpio6_0_analog_sel,
	output wire	gpio6_0_hys_trim,
	output wire	gpio6_0_hld_ovr,
	input wire	gpio6_0_in_h,
	output wire	gpio6_0_enable_h,
	input wire	gpio6_0_in,
	output wire	gpio6_0_hld_h_n,
	output wire	gpio6_0_enable_vdda_h,
	output wire	gpio6_0_analog_en,
	output wire	gpio6_0_enable_inp_h,
	output wire	gpio6_0_enable_vswitch_h,
	inout wire	gpio6_0_pad_a_noesd_h,
	inout wire	gpio6_0_pad_a_esd_0_h,
	inout wire	gpio6_0_pad_a_esd_1_h,
	input wire	gpio6_0_zero,
	input wire	gpio6_0_one,
	input wire	gpio6_1_tie_hi_esd,
	output wire	[2:0]	gpio6_1_dm,
	output wire	gpio6_1_slow,
	output wire	gpio6_1_oe_n,
	input wire	gpio6_1_tie_lo_esd,
	output wire	gpio6_1_inp_dis,
	output wire	gpio6_1_enable_vddio,
	output wire	gpio6_1_vtrip_sel,
	output wire	[1:0]	gpio6_1_ib_mode_sel,
	output wire	gpio6_1_out,
	output wire	[1:0]	gpio6_1_slew_ctl,
	output wire	gpio6_1_analog_pol,
	output wire	gpio6_1_analog_sel,
	output wire	gpio6_1_hys_trim,
	output wire	gpio6_1_hld_ovr,
	input wire	gpio6_1_in_h,
	output wire	gpio6_1_enable_h,
	input wire	gpio6_1_in,
	output wire	gpio6_1_hld_h_n,
	output wire	gpio6_1_enable_vdda_h,
	output wire	gpio6_1_analog_en,
	output wire	gpio6_1_enable_inp_h,
	output wire	gpio6_1_enable_vswitch_h,
	inout wire	gpio6_1_pad_a_noesd_h,
	inout wire	gpio6_1_pad_a_esd_0_h,
	inout wire	gpio6_1_pad_a_esd_1_h,
	input wire	gpio6_1_zero,
	input wire	gpio6_1_one,
	input wire	gpio6_2_tie_hi_esd,
	output wire	[2:0]	gpio6_2_dm,
	output wire	gpio6_2_slow,
	output wire	gpio6_2_oe_n,
	input wire	gpio6_2_tie_lo_esd,
	output wire	gpio6_2_inp_dis,
	output wire	gpio6_2_enable_vddio,
	output wire	gpio6_2_vtrip_sel,
	output wire	[1:0]	gpio6_2_ib_mode_sel,
	output wire	gpio6_2_out,
	output wire	[1:0]	gpio6_2_slew_ctl,
	output wire	gpio6_2_analog_pol,
	output wire	gpio6_2_analog_sel,
	output wire	gpio6_2_hys_trim,
	output wire	gpio6_2_hld_ovr,
	input wire	gpio6_2_in_h,
	output wire	gpio6_2_enable_h,
	input wire	gpio6_2_in,
	output wire	gpio6_2_hld_h_n,
	output wire	gpio6_2_enable_vdda_h,
	output wire	gpio6_2_analog_en,
	output wire	gpio6_2_enable_inp_h,
	output wire	gpio6_2_enable_vswitch_h,
	inout wire	gpio6_2_pad_a_noesd_h,
	inout wire	gpio6_2_pad_a_esd_0_h,
	inout wire	gpio6_2_pad_a_esd_1_h,
	input wire	gpio6_2_zero,
	input wire	gpio6_2_one,
	input wire	gpio6_3_tie_hi_esd,
	output wire	[2:0]	gpio6_3_dm,
	output wire	gpio6_3_slow,
	output wire	gpio6_3_oe_n,
	input wire	gpio6_3_tie_lo_esd,
	output wire	gpio6_3_inp_dis,
	output wire	gpio6_3_enable_vddio,
	output wire	gpio6_3_vtrip_sel,
	output wire	[1:0]	gpio6_3_ib_mode_sel,
	output wire	gpio6_3_out,
	output wire	[1:0]	gpio6_3_slew_ctl,
	output wire	gpio6_3_analog_pol,
	output wire	gpio6_3_analog_sel,
	output wire	gpio6_3_hys_trim,
	output wire	gpio6_3_hld_ovr,
	input wire	gpio6_3_in_h,
	output wire	gpio6_3_enable_h,
	input wire	gpio6_3_in,
	output wire	gpio6_3_hld_h_n,
	output wire	gpio6_3_enable_vdda_h,
	output wire	gpio6_3_analog_en,
	output wire	gpio6_3_enable_inp_h,
	output wire	gpio6_3_enable_vswitch_h,
	inout wire	gpio6_3_pad_a_noesd_h,
	inout wire	gpio6_3_pad_a_esd_0_h,
	inout wire	gpio6_3_pad_a_esd_1_h,
	input wire	gpio6_3_zero,
	input wire	gpio6_3_one,
	output wire	[4:0]	vref_w_ref_sel,
	inout wire	vref_w_vinref,
	output wire	vref_w_enable_h,
	output wire	vref_w_hld_h_n,
	output wire	vref_w_vrefgen_en,
	input wire	gpio6_4_tie_hi_esd,
	output wire	[2:0]	gpio6_4_dm,
	output wire	gpio6_4_slow,
	output wire	gpio6_4_oe_n,
	input wire	gpio6_4_tie_lo_esd,
	output wire	gpio6_4_inp_dis,
	output wire	gpio6_4_enable_vddio,
	output wire	gpio6_4_vtrip_sel,
	output wire	[1:0]	gpio6_4_ib_mode_sel,
	output wire	gpio6_4_out,
	output wire	[1:0]	gpio6_4_slew_ctl,
	output wire	gpio6_4_analog_pol,
	output wire	gpio6_4_analog_sel,
	output wire	gpio6_4_hys_trim,
	output wire	gpio6_4_hld_ovr,
	input wire	gpio6_4_in_h,
	output wire	gpio6_4_enable_h,
	input wire	gpio6_4_in,
	output wire	gpio6_4_hld_h_n,
	output wire	gpio6_4_enable_vdda_h,
	output wire	gpio6_4_analog_en,
	output wire	gpio6_4_enable_inp_h,
	output wire	gpio6_4_enable_vswitch_h,
	inout wire	gpio6_4_pad_a_noesd_h,
	inout wire	gpio6_4_pad_a_esd_0_h,
	inout wire	gpio6_4_pad_a_esd_1_h,
	input wire	gpio6_4_zero,
	input wire	gpio6_4_one,
	input wire	gpio6_5_tie_hi_esd,
	output wire	[2:0]	gpio6_5_dm,
	output wire	gpio6_5_slow,
	output wire	gpio6_5_oe_n,
	input wire	gpio6_5_tie_lo_esd,
	output wire	gpio6_5_inp_dis,
	output wire	gpio6_5_enable_vddio,
	output wire	gpio6_5_vtrip_sel,
	output wire	[1:0]	gpio6_5_ib_mode_sel,
	output wire	gpio6_5_out,
	output wire	[1:0]	gpio6_5_slew_ctl,
	output wire	gpio6_5_analog_pol,
	output wire	gpio6_5_analog_sel,
	output wire	gpio6_5_hys_trim,
	output wire	gpio6_5_hld_ovr,
	input wire	gpio6_5_in_h,
	output wire	gpio6_5_enable_h,
	input wire	gpio6_5_in,
	output wire	gpio6_5_hld_h_n,
	output wire	gpio6_5_enable_vdda_h,
	output wire	gpio6_5_analog_en,
	output wire	gpio6_5_enable_inp_h,
	output wire	gpio6_5_enable_vswitch_h,
	inout wire	gpio6_5_pad_a_noesd_h,
	inout wire	gpio6_5_pad_a_esd_0_h,
	inout wire	gpio6_5_pad_a_esd_1_h,
	input wire	gpio6_5_zero,
	input wire	gpio6_5_one,
	input wire	gpio6_6_tie_hi_esd,
	output wire	[2:0]	gpio6_6_dm,
	output wire	gpio6_6_slow,
	output wire	gpio6_6_oe_n,
	input wire	gpio6_6_tie_lo_esd,
	output wire	gpio6_6_inp_dis,
	output wire	gpio6_6_enable_vddio,
	output wire	gpio6_6_vtrip_sel,
	output wire	[1:0]	gpio6_6_ib_mode_sel,
	output wire	gpio6_6_out,
	output wire	[1:0]	gpio6_6_slew_ctl,
	output wire	gpio6_6_analog_pol,
	output wire	gpio6_6_analog_sel,
	output wire	gpio6_6_hys_trim,
	output wire	gpio6_6_hld_ovr,
	input wire	gpio6_6_in_h,
	output wire	gpio6_6_enable_h,
	input wire	gpio6_6_in,
	output wire	gpio6_6_hld_h_n,
	output wire	gpio6_6_enable_vdda_h,
	output wire	gpio6_6_analog_en,
	output wire	gpio6_6_enable_inp_h,
	output wire	gpio6_6_enable_vswitch_h,
	inout wire	gpio6_6_pad_a_noesd_h,
	inout wire	gpio6_6_pad_a_esd_0_h,
	inout wire	gpio6_6_pad_a_esd_1_h,
	input wire	gpio6_6_zero,
	input wire	gpio6_6_one,
	input wire	gpio6_7_tie_hi_esd,
	output wire	[2:0]	gpio6_7_dm,
	output wire	gpio6_7_slow,
	output wire	gpio6_7_oe_n,
	input wire	gpio6_7_tie_lo_esd,
	output wire	gpio6_7_inp_dis,
	output wire	gpio6_7_enable_vddio,
	output wire	gpio6_7_vtrip_sel,
	output wire	[1:0]	gpio6_7_ib_mode_sel,
	output wire	gpio6_7_out,
	output wire	[1:0]	gpio6_7_slew_ctl,
	output wire	gpio6_7_analog_pol,
	output wire	gpio6_7_analog_sel,
	output wire	gpio6_7_hys_trim,
	output wire	gpio6_7_hld_ovr,
	input wire	gpio6_7_in_h,
	output wire	gpio6_7_enable_h,
	input wire	gpio6_7_in,
	output wire	gpio6_7_hld_h_n,
	output wire	gpio6_7_enable_vdda_h,
	output wire	gpio6_7_analog_en,
	output wire	gpio6_7_enable_inp_h,
	output wire	gpio6_7_enable_vswitch_h,
	inout wire	gpio6_7_pad_a_noesd_h,
	inout wire	gpio6_7_pad_a_esd_0_h,
	inout wire	gpio6_7_pad_a_esd_1_h,
	input wire	gpio6_7_zero,
	input wire	gpio6_7_one,
	input wire	gpio7_0_tie_lo_esd,
	input wire	gpio7_0_in,
	input wire	gpio7_0_tie_hi_esd,
	output wire	gpio7_0_enable_vddio,
	output wire	gpio7_0_slow,
	inout wire	gpio7_0_pad_a_esd_0_h,
	inout wire	gpio7_0_pad_a_esd_1_h,
	inout wire	gpio7_0_pad_a_noesd_h,
	output wire	gpio7_0_analog_en,
	output wire	gpio7_0_analog_pol,
	output wire	gpio7_0_inp_dis,
	output wire	gpio7_0_enable_inp_h,
	output wire	gpio7_0_enable_h,
	output wire	gpio7_0_hld_h_n,
	output wire	gpio7_0_analog_sel,
	output wire	[2:0]	gpio7_0_dm,
	output wire	gpio7_0_hld_ovr,
	output wire	gpio7_0_out,
	output wire	gpio7_0_enable_vswitch_h,
	output wire	gpio7_0_enable_vdda_h,
	output wire	gpio7_0_vtrip_sel,
	output wire	gpio7_0_ib_mode_sel,
	output wire	gpio7_0_oe_n,
	input wire	gpio7_0_in_h,
	input wire	gpio7_0_zero,
	input wire	gpio7_0_one,
	input wire	gpio7_1_tie_lo_esd,
	input wire	gpio7_1_in,
	input wire	gpio7_1_tie_hi_esd,
	output wire	gpio7_1_enable_vddio,
	output wire	gpio7_1_slow,
	inout wire	gpio7_1_pad_a_esd_0_h,
	inout wire	gpio7_1_pad_a_esd_1_h,
	inout wire	gpio7_1_pad_a_noesd_h,
	output wire	gpio7_1_analog_en,
	output wire	gpio7_1_analog_pol,
	output wire	gpio7_1_inp_dis,
	output wire	gpio7_1_enable_inp_h,
	output wire	gpio7_1_enable_h,
	output wire	gpio7_1_hld_h_n,
	output wire	gpio7_1_analog_sel,
	output wire	[2:0]	gpio7_1_dm,
	output wire	gpio7_1_hld_ovr,
	output wire	gpio7_1_out,
	output wire	gpio7_1_enable_vswitch_h,
	output wire	gpio7_1_enable_vdda_h,
	output wire	gpio7_1_vtrip_sel,
	output wire	gpio7_1_ib_mode_sel,
	output wire	gpio7_1_oe_n,
	input wire	gpio7_1_in_h,
	input wire	gpio7_1_zero,
	input wire	gpio7_1_one,
	input wire	gpio7_2_tie_lo_esd,
	input wire	gpio7_2_in,
	input wire	gpio7_2_tie_hi_esd,
	output wire	gpio7_2_enable_vddio,
	output wire	gpio7_2_slow,
	inout wire	gpio7_2_pad_a_esd_0_h,
	inout wire	gpio7_2_pad_a_esd_1_h,
	inout wire	gpio7_2_pad_a_noesd_h,
	output wire	gpio7_2_analog_en,
	output wire	gpio7_2_analog_pol,
	output wire	gpio7_2_inp_dis,
	output wire	gpio7_2_enable_inp_h,
	output wire	gpio7_2_enable_h,
	output wire	gpio7_2_hld_h_n,
	output wire	gpio7_2_analog_sel,
	output wire	[2:0]	gpio7_2_dm,
	output wire	gpio7_2_hld_ovr,
	output wire	gpio7_2_out,
	output wire	gpio7_2_enable_vswitch_h,
	output wire	gpio7_2_enable_vdda_h,
	output wire	gpio7_2_vtrip_sel,
	output wire	gpio7_2_ib_mode_sel,
	output wire	gpio7_2_oe_n,
	input wire	gpio7_2_in_h,
	input wire	gpio7_2_zero,
	input wire	gpio7_2_one,
	input wire	gpio7_3_tie_lo_esd,
	input wire	gpio7_3_in,
	input wire	gpio7_3_tie_hi_esd,
	output wire	gpio7_3_enable_vddio,
	output wire	gpio7_3_slow,
	inout wire	gpio7_3_pad_a_esd_0_h,
	inout wire	gpio7_3_pad_a_esd_1_h,
	inout wire	gpio7_3_pad_a_noesd_h,
	output wire	gpio7_3_analog_en,
	output wire	gpio7_3_analog_pol,
	output wire	gpio7_3_inp_dis,
	output wire	gpio7_3_enable_inp_h,
	output wire	gpio7_3_enable_h,
	output wire	gpio7_3_hld_h_n,
	output wire	gpio7_3_analog_sel,
	output wire	[2:0]	gpio7_3_dm,
	output wire	gpio7_3_hld_ovr,
	output wire	gpio7_3_out,
	output wire	gpio7_3_enable_vswitch_h,
	output wire	gpio7_3_enable_vdda_h,
	output wire	gpio7_3_vtrip_sel,
	output wire	gpio7_3_ib_mode_sel,
	output wire	gpio7_3_oe_n,
	input wire	gpio7_3_in_h,
	input wire	gpio7_3_zero,
	input wire	gpio7_3_one,
	input wire	gpio7_4_tie_lo_esd,
	input wire	gpio7_4_in,
	input wire	gpio7_4_tie_hi_esd,
	output wire	gpio7_4_enable_vddio,
	output wire	gpio7_4_slow,
	inout wire	gpio7_4_pad_a_esd_0_h,
	inout wire	gpio7_4_pad_a_esd_1_h,
	inout wire	gpio7_4_pad_a_noesd_h,
	output wire	gpio7_4_analog_en,
	output wire	gpio7_4_analog_pol,
	output wire	gpio7_4_inp_dis,
	output wire	gpio7_4_enable_inp_h,
	output wire	gpio7_4_enable_h,
	output wire	gpio7_4_hld_h_n,
	output wire	gpio7_4_analog_sel,
	output wire	[2:0]	gpio7_4_dm,
	output wire	gpio7_4_hld_ovr,
	output wire	gpio7_4_out,
	output wire	gpio7_4_enable_vswitch_h,
	output wire	gpio7_4_enable_vdda_h,
	output wire	gpio7_4_vtrip_sel,
	output wire	gpio7_4_ib_mode_sel,
	output wire	gpio7_4_oe_n,
	input wire	gpio7_4_in_h,
	input wire	gpio7_4_zero,
	input wire	gpio7_4_one,
	input wire	gpio7_5_tie_lo_esd,
	input wire	gpio7_5_in,
	input wire	gpio7_5_tie_hi_esd,
	output wire	gpio7_5_enable_vddio,
	output wire	gpio7_5_slow,
	inout wire	gpio7_5_pad_a_esd_0_h,
	inout wire	gpio7_5_pad_a_esd_1_h,
	inout wire	gpio7_5_pad_a_noesd_h,
	output wire	gpio7_5_analog_en,
	output wire	gpio7_5_analog_pol,
	output wire	gpio7_5_inp_dis,
	output wire	gpio7_5_enable_inp_h,
	output wire	gpio7_5_enable_h,
	output wire	gpio7_5_hld_h_n,
	output wire	gpio7_5_analog_sel,
	output wire	[2:0]	gpio7_5_dm,
	output wire	gpio7_5_hld_ovr,
	output wire	gpio7_5_out,
	output wire	gpio7_5_enable_vswitch_h,
	output wire	gpio7_5_enable_vdda_h,
	output wire	gpio7_5_vtrip_sel,
	output wire	gpio7_5_ib_mode_sel,
	output wire	gpio7_5_oe_n,
	input wire	gpio7_5_in_h,
	input wire	gpio7_5_zero,
	input wire	gpio7_5_one,
	input wire	gpio7_6_tie_lo_esd,
	input wire	gpio7_6_in,
	input wire	gpio7_6_tie_hi_esd,
	output wire	gpio7_6_enable_vddio,
	output wire	gpio7_6_slow,
	inout wire	gpio7_6_pad_a_esd_0_h,
	inout wire	gpio7_6_pad_a_esd_1_h,
	inout wire	gpio7_6_pad_a_noesd_h,
	output wire	gpio7_6_analog_en,
	output wire	gpio7_6_analog_pol,
	output wire	gpio7_6_inp_dis,
	output wire	gpio7_6_enable_inp_h,
	output wire	gpio7_6_enable_h,
	output wire	gpio7_6_hld_h_n,
	output wire	gpio7_6_analog_sel,
	output wire	[2:0]	gpio7_6_dm,
	output wire	gpio7_6_hld_ovr,
	output wire	gpio7_6_out,
	output wire	gpio7_6_enable_vswitch_h,
	output wire	gpio7_6_enable_vdda_h,
	output wire	gpio7_6_vtrip_sel,
	output wire	gpio7_6_ib_mode_sel,
	output wire	gpio7_6_oe_n,
	input wire	gpio7_6_in_h,
	input wire	gpio7_6_zero,
	input wire	gpio7_6_one,
	input wire	gpio7_7_tie_lo_esd,
	input wire	gpio7_7_in,
	input wire	gpio7_7_tie_hi_esd,
	output wire	gpio7_7_enable_vddio,
	output wire	gpio7_7_slow,
	inout wire	gpio7_7_pad_a_esd_0_h,
	inout wire	gpio7_7_pad_a_esd_1_h,
	inout wire	gpio7_7_pad_a_noesd_h,
	output wire	gpio7_7_analog_en,
	output wire	gpio7_7_analog_pol,
	output wire	gpio7_7_inp_dis,
	output wire	gpio7_7_enable_inp_h,
	output wire	gpio7_7_enable_h,
	output wire	gpio7_7_hld_h_n,
	output wire	gpio7_7_analog_sel,
	output wire	[2:0]	gpio7_7_dm,
	output wire	gpio7_7_hld_ovr,
	output wire	gpio7_7_out,
	output wire	gpio7_7_enable_vswitch_h,
	output wire	gpio7_7_enable_vdda_h,
	output wire	gpio7_7_vtrip_sel,
	output wire	gpio7_7_ib_mode_sel,
	output wire	gpio7_7_oe_n,
	input wire	gpio7_7_in_h,
	input wire	gpio7_7_zero,
	input wire	gpio7_7_one,
	output wire	muxsplit_sw_hld_vdda_h_n,
	output wire	muxsplit_sw_enable_vdda_h,
	output wire	muxsplit_sw_switch_aa_sl,
	output wire	muxsplit_sw_switch_aa_s0,
	output wire	muxsplit_sw_switch_bb_s0,
	output wire	muxsplit_sw_switch_bb_sl,
	output wire	muxsplit_sw_switch_bb_sr,
	output wire	muxsplit_sw_switch_aa_sr
);

    wire xclk;
    
    // Sync reset
    reg [1:0] xrst_n_d;
    wire xrst_n;
    always @(posedge xclk) begin
        xrst_n_d <= {xrst_n_d[0], resetb_xres_n};
    end
    assign xrst_n = xrst_n_d[1];
    
    //wire xrst_n;
    //assign xrst_n = resetb_xres_n;
    
    (* dont_touch *) wire porb_h;
    
    sky130_ef_ip__simple_por4x simple_por4x (
    `ifdef FUNCTIONAL
    `ifdef USE_POWER_PINS
        .vdd3v3 (DVPWR),
        .vdd1v8 (AVPWR),
        .vss3v3 (DVGND),
        .vss1v8 (AVGND),
    `endif
    `endif
        .porb_h (porb_h),
        .porb_l (),
        .por_l  ()
    );
    
    parameter FABRIC_NUM_IO_WEST = 64;
    
    wire [FABRIC_NUM_IO_WEST-1:0] fabric_io_in;
    wire [FABRIC_NUM_IO_WEST-1:0] fabric_io_out;
    wire [FABRIC_NUM_IO_WEST-1:0] fabric_io_oe;

    wire [FABRIC_NUM_IO_WEST-1:0] fabric_io_config_bit0;
    wire [FABRIC_NUM_IO_WEST-1:0] fabric_io_config_bit1;
    wire [FABRIC_NUM_IO_WEST-1:0] fabric_io_config_bit2;
    wire [FABRIC_NUM_IO_WEST-1:0] fabric_io_config_bit3;

    wire fpga_mode_i;
    wire config_busy_o;

    wire fpga_sclk_in;
    wire fpga_sclk_out;
    wire fpga_sclk_oe, fpga_sclk_oeb;
    assign fpga_sclk_oeb = !fpga_sclk_oe;
    
    wire fpga_cs_n_in;
    wire fpga_cs_n_out;
    wire fpga_cs_n_oe, fpga_cs_n_oeb;
    assign fpga_cs_n_oeb = !fpga_cs_n_oe;
    
    wire fpga_mosi_in;
    wire fpga_mosi_out;
    wire fpga_mosi_oe, fpga_mosi_oeb;
    assign fpga_mosi_oeb = !fpga_mosi_oe;
    
    wire fpga_miso_in;
    wire fpga_miso_out;
    wire fpga_miso_oe, fpga_miso_oeb;
    assign fpga_miso_oeb = !fpga_miso_oe;
    
    // ADC 0
    wire        fabric_adc0_cmp_i;
    wire        fabric_adc0_hold_o;
    wire        fabric_adc0_reset_o;
    wire [11:0] fabric_adc0_value_o;

    // ADC 1
    wire        fabric_adc1_cmp_i;
    wire        fabric_adc1_hold_o;
    wire        fabric_adc1_reset_o;
    wire [11:0] fabric_adc1_value_o;

    // DAC 0
    wire [7:0]  fabric_dac0_value_o;
    wire        fabric_dac0_enable_o;

    // DAC 1
    wire [7:0]  fabric_dac1_value_o;
    wire        fabric_dac1_enable_o;

    panamax_fpga_core #(
        .FABRIC_NUM_IO_WEST (FABRIC_NUM_IO_WEST)
    ) panamax_fpga_core (
    `ifdef USE_POWER_PINS
        .VPWR   (DVPWR),
        .VGND   (DVGND),
    `endif
    
        .clk_i      (xclk),
        .rst_ni     (xrst_n),
        
        // FPGA config
        .fpga_sclk_i        (fpga_sclk_in),
        .fpga_sclk_o        (fpga_sclk_out),
        .fpga_sclk_oe_o     (fpga_sclk_oe),

        .fpga_cs_n_i        (fpga_cs_n_in),
        .fpga_cs_n_o        (fpga_cs_n_out),
        .fpga_cs_n_oe_o     (fpga_cs_n_oe),

        .fpga_mosi_i        (fpga_mosi_in),
        .fpga_mosi_o        (fpga_mosi_out),
        .fpga_mosi_oe_o     (fpga_mosi_oe),

        .fpga_miso_i        (fpga_miso_in),
        .fpga_miso_o        (fpga_miso_out),
        .fpga_miso_oe_o     (fpga_miso_oe),
        
        // FPGA config mode
        // if mode == 0: SPI controller
        // if mode == 1: SPI receiver
        .fpga_mode_i,
        .config_busy_o,
        
        // ADC 0
        .fabric_adc0_cmp_i      (fabric_adc0_cmp_i),
        .fabric_adc0_hold_o     (fabric_adc0_hold_o),
        .fabric_adc0_reset_o    (fabric_adc0_reset_o),
        .fabric_adc0_value_o    (fabric_adc0_value_o),

        // ADC 1
        .fabric_adc1_cmp_i      (fabric_adc1_cmp_i),
        .fabric_adc1_hold_o     (fabric_adc1_hold_o),
        .fabric_adc1_reset_o    (fabric_adc1_reset_o),
        .fabric_adc1_value_o    (fabric_adc1_value_o),

        // DAC 0
        .fabric_dac0_value_o    (fabric_dac0_value_o),
        .fabric_dac0_enable_o   (fabric_dac0_enable_o),

        // DAC 1
        .fabric_dac1_value_o    (fabric_dac1_value_o),
        .fabric_dac1_enable_o   (fabric_dac1_enable_o),

        // Fabric I/O
        .fabric_io_in_i     (fabric_io_in),
        .fabric_io_out_o    (fabric_io_out),
        .fabric_io_oe_o     (fabric_io_oe),
        
        .fabric_io_config_bit0_o    (fabric_io_config_bit0),
        .fabric_io_config_bit1_o    (fabric_io_config_bit1),
        .fabric_io_config_bit2_o    (fabric_io_config_bit2),
        .fabric_io_config_bit3_o    (fabric_io_config_bit3)
    );

    (* keep *) sky130_ef_ip__rdac3v_8bit dac0 (
    /*`ifdef USE_POWER_PINS
        .vdd    (AVPWR),
        .vss    (AVGND),
        .dvdd   (DVPWR),
        .dvss   (DVGND),

        .Vhigh  (AVPWR),
        .Vlow   (AVGND),

        .out    (xi1_core),
    `endif*/

       .b   (fabric_dac0_value_o),
       .ena (fabric_dac0_enable_o)
    );
    
    (* keep *) sky130_ef_ip__rdac3v_8bit dac1 (
    /*`ifdef USE_POWER_PINS
        .vdd    (AVPWR),
        .vss    (AVGND),
        .dvdd   (DVPWR),
        .dvss   (DVGND),

        .Vhigh  (AVPWR),
        .Vlow   (AVGND),

        .out    (xo1_core),
    `endif*/

       .b   (fabric_dac1_value_o),
       .ena (fabric_dac1_enable_o)
    );
    
    `ifdef USE_POWER_PINS
    wire adc0_vref;
    wire adc1_vref;
    `endif
    
    (* keep *) res_div res_div0 (
    `ifdef USE_POWER_PINS
        .vdda  (AVPWR),
        .vssa  (AVGND),
        .vref  (adc0_vref)
    `endif
    );
    
    (* keep *) res_div res_div1 (
    `ifdef USE_POWER_PINS
        .vdda  (AVPWR),
        .vssa  (AVGND),
        .vref  (adc1_vref)
    `endif
    );
    
    (* keep *) sky130_ef_ip__adc3v_12bit adc0 (
    `ifdef USE_POWER_PINS
        .vccd0  (DVPWR),
        .vssd0  (DVGND),
        .vdda0  (AVPWR),
        .vssa0  (AVGND),
       
        .adc_trim   (AVGND),
        .adc_vCM    (adc0_vref),
        .adc_vrefL  (AVGND),
        .adc_vrefH  (AVPWR),
        .adc_in     (xi0_core),
    `endif

       .adc_ena        (1'b1),
       .adc_reset      (fabric_adc0_reset_o),
       .adc_hold       (fabric_adc0_hold_o),
       .adc_dac_val    (fabric_adc0_value_o),
       .adc_comp_out   (fabric_adc0_cmp_i)
    );
    
    (* keep *) sky130_ef_ip__adc3v_12bit adc1 (
    `ifdef USE_POWER_PINS
        .vccd0  (DVPWR),
        .vssd0  (DVGND),
        .vdda0  (AVPWR),
        .vssa0  (AVGND),
       
        .adc_trim   (AVGND),
        .adc_vCM    (adc1_vref),
        .adc_vrefL  (AVGND),
        .adc_vrefH  (AVPWR),
        .adc_in     (xo0_core),
    `endif

       .adc_ena        (1'b1),
       .adc_reset      (fabric_adc1_reset_o),
       .adc_hold       (fabric_adc1_hold_o),
       .adc_dac_val    (fabric_adc1_value_o),
       .adc_comp_out   (fabric_adc1_cmp_i)
    );
    
    wire [0:0] unused;

    `include "gpio_mapping.v"
    
    // GPIO mapping for SIO 0 & 1

    // SIO 0 (GPIO 72)
    //assign TODO       = sio_in[0];
    assign sio_out[0]           = gpio0_0_zero;
    assign sio_oe_n[0]          = gpio0_0_one;
    assign sio_inp_dis[0]       = gpio0_0_one;
    assign sio_vtrip_sel[0]     = gpio0_0_zero;
    assign sio_slow[0]          = gpio0_0_zero;
    assign sio_hld_ovr[0]       = gpio0_0_zero;
    assign sio_dm0              = {gpio0_0_one, gpio0_0_one, gpio0_0_zero};
    // assign sio_enable_vddio[0]  = 1'b1; // Not exported from panamax
    // assign sio_enable_inp_h[0]  = sio_tie_lo_esd[0]; // Not exported from panamax
    assign sio_enable_h         = porb_h;
    assign sio_hld_h_n[0]       = gpio0_0_tie_hi_esd;
    assign sio_enable_vdda_h    = porb_h;
    assign sio_ibuf_sel[0]      = gpio0_0_zero;
    assign sio_vreg_en[0]       = gpio0_0_zero; // TODO

    assign sio_hld_h_n_refgen   = gpio0_0_tie_hi_esd; 
    assign sio_ibuf_sel_refgen  = gpio0_0_zero; // TODO
    assign sio_vtrip_sel_refgen = gpio0_0_zero; // TODO
    assign sio_dft_refgen       = gpio0_0_zero; // disable ADFT
    // assign sio_vohref           = 1'b1; // TODO: Analog connection -> ground to vssa
    // sio_vinref_dft // ADFT test point -> floating
    // voutref_dft // ADFT test point -> our reference for vcm


    // SIO 1 (GPIO 73)
    //assign TODO           = sio_in[1];
    assign sio_out[1]               = gpio0_0_zero;
    assign sio_oe_n[1]              = gpio0_0_one;
    assign sio_inp_dis[1]           = gpio0_0_one;
    assign sio_vtrip_sel[1]         = gpio0_0_zero;
    assign sio_slow[1]              = gpio0_0_zero;
    assign sio_hld_ovr[1]           = gpio0_0_zero;
    assign sio_dm1                  = {gpio0_0_one, gpio0_0_one, gpio0_0_zero};
    // assign sio_enable_vddio[1]      = 1'b1; // Not exported from panamax
    // assign sio_enable_inp_h[1]      = sio_tie_lo_esd[1]; // Not exported from panamax
    assign sio_hld_h_n[1]           = gpio0_0_tie_hi_esd;
    assign sio_ibuf_sel[1]          = gpio0_0_zero;
    assign sio_vreg_en[1]           = gpio0_0_zero; // TODO
    
    assign sio_voh_sel              = {gpio0_0_one, gpio0_0_zero, gpio0_0_zero}; // n = Rtap/Rtotal = 1
    assign sio_vref_sel             = {gpio0_0_zero, gpio0_0_zero}; // Vohref
    assign sio_vreg_en_refgen       = gpio0_0_zero; // disable refgen
    

    // resetb PAD
    wire xres_loop;
    wire xres_vss_loop;
    assign xres_loop = resetb_tie_weak_hi_h;
    assign xres_loop = resetb_pad_a_esd_h;
    assign resetb_disable_pullup_h = xres_vss_loop;
    // assign resetb_tie_hi_esd =
    assign xres_vss_loop = resetb_tie_lo_esd;
    assign resetb_inp_sel_h = xres_vss_loop;
    assign resetb_en_vddio_sig_h = xres_vss_loop;
    assign resetb_filt_in_h = xres_vss_loop;
    assign resetb_pullup_h = xres_vss_loop;
    assign resetb_enable_h = porb_h ;
    assign resetb_enable_vddio = select_one;

    // muxsplit
    assign muxsplit_ne_enable_vdda_h = porb_h ;
    assign muxsplit_ne_hld_vdda_h_n = gpio2_7_tie_hi_esd; // nearest tie hi esd
    assign muxsplit_nw_enable_vdda_h = porb_h ;
    assign muxsplit_nw_hld_vdda_h_n = gpio5_0_tie_hi_esd; // nearest tie hi esd
    assign muxsplit_se_enable_vdda_h = porb_h ;
    assign muxsplit_se_hld_vdda_h_n = gpio0_0_tie_hi_esd; // nearest tie hi esd
    assign muxsplit_sw_enable_vdda_h = porb_h ;
    assign muxsplit_sw_hld_vdda_h_n = gpio7_7_tie_hi_esd; // nearest tie hi esd

    // Can be used to route analog signals in the padring
    assign muxsplit_ne_switch_aa_sl = 1'b0;
    assign muxsplit_ne_switch_aa_s0 = 1'b0;
    assign muxsplit_ne_switch_bb_s0 = 1'b0;
    assign muxsplit_ne_switch_bb_sl = 1'b0;
    assign muxsplit_ne_switch_bb_sr = 1'b0;
    assign muxsplit_ne_switch_aa_sr = 1'b0;

    assign muxsplit_nw_switch_aa_sl = 1'b0;
    assign muxsplit_nw_switch_aa_s0 = 1'b0;
    assign muxsplit_nw_switch_bb_s0 = 1'b0;
    assign muxsplit_nw_switch_bb_sl = 1'b0;
    assign muxsplit_nw_switch_bb_sr = 1'b0;
    assign muxsplit_nw_switch_aa_sr = 1'b0;

    assign muxsplit_se_switch_aa_sl = 1'b0;
    assign muxsplit_se_switch_aa_s0 = 1'b0;
    assign muxsplit_se_switch_bb_s0 = 1'b0;
    assign muxsplit_se_switch_bb_sl = 1'b0;
    assign muxsplit_se_switch_bb_sr = 1'b0;
    assign muxsplit_se_switch_aa_sr = 1'b0;

    assign muxsplit_sw_switch_aa_sl = 1'b0;
    assign muxsplit_sw_switch_aa_s0 = 1'b0;
    assign muxsplit_sw_switch_bb_s0 = 1'b0;
    assign muxsplit_sw_switch_bb_sl = 1'b0;
    assign muxsplit_sw_switch_bb_sr = 1'b0;
    assign muxsplit_sw_switch_aa_sr = 1'b0;

    // vrefs
    assign vref_e_enable_h = porb_h;
    assign vref_e_hld_h_n = gpio1_4_tie_hi_esd; // nearest tie hi esd
    assign vref_w_enable_h = porb_h;
    assign vref_w_hld_h_n = gpio6_4_tie_hi_esd; // nearest tie hi esd

    // Doesn't matter, we don't use vrefs
    assign vref_e_ref_sel = 5'b01111;
    assign vref_e_vrefgen_en = 1'b1;

    assign vref_w_ref_sel = 5'b01111;
    assign vref_w_vrefgen_en = 1'b1;
    
    // analog vref_e_vinref
    // analog vref_w_vinref

    // Select
    //assign mgmt_select = select_in;
    assign select_enable_vddio      = select_one;
    assign select_slow              = select_zero;
    assign select_analog_en         = select_zero;
    assign select_analog_pol        = select_zero;
    assign select_inp_dis           = select_zero;
    assign select_enable_inp_h      = select_tie_lo_esd;
    assign select_enable_h          = porb_h;
    assign select_hld_h_n           = select_tie_hi_esd;
    assign select_analog_sel        = select_zero;
    assign select_dm                = {select_zero, select_one, select_one};
    assign select_hld_ovr           = select_zero;
    assign select_out               = select_zero;
    assign select_enable_vswitch_h  = select_tie_hi_esd;
    assign select_enable_vdda_h     = porb_h;
    assign select_vtrip_sel         = select_zero;
    assign select_ib_mode_sel       = select_zero;
    assign select_oe_n              = select_zero;
    
    // Power detector is not used
    assign pwrdet_in1_vddio_hv = 1'b0;
    assign pwrdet_in2_vddd_hv = 1'b0;
    assign pwrdet_in1_vddd_hv = 1'b0;
    assign pwrdet_in3_vddd_hv = 1'b0;
    assign pwrdet_in2_vddio_hv = 1'b0;
    assign pwrdet_in3_vddio_hv = 1'b0;
    assign pwrdet_rst_por_hv_n = 1'b0;
    
    (* keep *) manual_routing manual_routing (
    /*`ifdef USE_POWER_PINS
        .DVPWR  (DVPWR),
        .DVGND  (DVGND)
    `endif*/
    );

endmodule

`default_nettype wire
