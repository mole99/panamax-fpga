module res_div (
    `ifdef USE_POWER_PINS
    inout vdda,
    inout vssa,
    inout vref
    `endif
);

endmodule
