module res_div (
    `ifdef USE_POWER_PINS
    inout vdda,
    inout vssa,
    inout vsub,
    inout vref
    `endif
);

endmodule
