VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO dll
  CLASS BLOCK ;
  FOREIGN dll ;
  ORIGIN 0.000 0.000 ;
  SIZE 135.000 BY 110.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 41.040 5.200 42.640 103.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 81.040 5.200 82.640 103.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 121.040 5.200 122.640 103.600 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 5.200 22.640 103.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 61.040 5.200 62.640 103.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 101.040 5.200 102.640 103.600 ;
    END
  END VPWR
  PIN clockp[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 5.480 4.000 6.080 ;
    END
  END clockp[0]
  PIN clockp[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 4.000 11.520 ;
    END
  END clockp[1]
  PIN dco
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.393000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 4.000 65.920 ;
    END
  END dco
  PIN div[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.360 4.000 16.960 ;
    END
  END div[0]
  PIN div[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.800 4.000 22.400 ;
    END
  END div[1]
  PIN div[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.621000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END div[2]
  PIN div[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.621000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 4.000 33.280 ;
    END
  END div[3]
  PIN div[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 4.000 38.720 ;
    END
  END div[4]
  PIN div[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 4.000 44.160 ;
    END
  END div[5]
  PIN div[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.000 4.000 49.600 ;
    END
  END div[6]
  PIN div[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.499500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END div[7]
  PIN enable
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.880 4.000 60.480 ;
    END
  END enable
  PIN ext_trim[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.760 4.000 71.360 ;
    END
  END ext_trim[0]
  PIN ext_trim[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 36.890 106.000 37.170 110.000 ;
    END
  END ext_trim[10]
  PIN ext_trim[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 47.010 106.000 47.290 110.000 ;
    END
  END ext_trim[11]
  PIN ext_trim[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 57.130 106.000 57.410 110.000 ;
    END
  END ext_trim[12]
  PIN ext_trim[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 67.250 106.000 67.530 110.000 ;
    END
  END ext_trim[13]
  PIN ext_trim[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 77.370 106.000 77.650 110.000 ;
    END
  END ext_trim[14]
  PIN ext_trim[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 87.490 106.000 87.770 110.000 ;
    END
  END ext_trim[15]
  PIN ext_trim[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 97.610 106.000 97.890 110.000 ;
    END
  END ext_trim[16]
  PIN ext_trim[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 107.730 106.000 108.010 110.000 ;
    END
  END ext_trim[17]
  PIN ext_trim[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 117.850 106.000 118.130 110.000 ;
    END
  END ext_trim[18]
  PIN ext_trim[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 127.970 106.000 128.250 110.000 ;
    END
  END ext_trim[19]
  PIN ext_trim[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.200 4.000 76.800 ;
    END
  END ext_trim[1]
  PIN ext_trim[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 131.000 97.960 135.000 98.560 ;
    END
  END ext_trim[20]
  PIN ext_trim[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 131.000 80.280 135.000 80.880 ;
    END
  END ext_trim[21]
  PIN ext_trim[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 131.000 62.600 135.000 63.200 ;
    END
  END ext_trim[22]
  PIN ext_trim[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 131.000 44.920 135.000 45.520 ;
    END
  END ext_trim[23]
  PIN ext_trim[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 131.000 27.240 135.000 27.840 ;
    END
  END ext_trim[24]
  PIN ext_trim[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 131.000 9.560 135.000 10.160 ;
    END
  END ext_trim[25]
  PIN ext_trim[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END ext_trim[2]
  PIN ext_trim[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.080 4.000 87.680 ;
    END
  END ext_trim[3]
  PIN ext_trim[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 4.000 93.120 ;
    END
  END ext_trim[4]
  PIN ext_trim[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.960 4.000 98.560 ;
    END
  END ext_trim[5]
  PIN ext_trim[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.400 4.000 104.000 ;
    END
  END ext_trim[6]
  PIN ext_trim[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 6.530 106.000 6.810 110.000 ;
    END
  END ext_trim[7]
  PIN ext_trim[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 16.650 106.000 16.930 110.000 ;
    END
  END ext_trim[8]
  PIN ext_trim[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 26.770 106.000 27.050 110.000 ;
    END
  END ext_trim[9]
  PIN osc
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 100.830 0.000 101.110 4.000 ;
    END
  END osc
  PIN resetb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 33.670 0.000 33.950 4.000 ;
    END
  END resetb
  OBS
      LAYER nwell ;
        RECT 5.330 5.355 129.450 103.445 ;
      LAYER li1 ;
        RECT 5.520 5.355 129.260 103.445 ;
      LAYER met1 ;
        RECT 0.990 5.200 132.410 106.720 ;
      LAYER met2 ;
        RECT 1.010 105.720 6.250 106.750 ;
        RECT 7.090 105.720 16.370 106.750 ;
        RECT 17.210 105.720 26.490 106.750 ;
        RECT 27.330 105.720 36.610 106.750 ;
        RECT 37.450 105.720 46.730 106.750 ;
        RECT 47.570 105.720 56.850 106.750 ;
        RECT 57.690 105.720 66.970 106.750 ;
        RECT 67.810 105.720 77.090 106.750 ;
        RECT 77.930 105.720 87.210 106.750 ;
        RECT 88.050 105.720 97.330 106.750 ;
        RECT 98.170 105.720 107.450 106.750 ;
        RECT 108.290 105.720 117.570 106.750 ;
        RECT 118.410 105.720 127.690 106.750 ;
        RECT 128.530 105.720 132.380 106.750 ;
        RECT 1.010 4.280 132.380 105.720 ;
        RECT 1.010 4.000 33.390 4.280 ;
        RECT 34.230 4.000 100.550 4.280 ;
        RECT 101.390 4.000 132.380 4.280 ;
      LAYER met3 ;
        RECT 4.400 103.000 131.000 103.865 ;
        RECT 0.985 98.960 131.000 103.000 ;
        RECT 4.400 97.560 130.600 98.960 ;
        RECT 0.985 93.520 131.000 97.560 ;
        RECT 4.400 92.120 131.000 93.520 ;
        RECT 0.985 88.080 131.000 92.120 ;
        RECT 4.400 86.680 131.000 88.080 ;
        RECT 0.985 82.640 131.000 86.680 ;
        RECT 4.400 81.280 131.000 82.640 ;
        RECT 4.400 81.240 130.600 81.280 ;
        RECT 0.985 79.880 130.600 81.240 ;
        RECT 0.985 77.200 131.000 79.880 ;
        RECT 4.400 75.800 131.000 77.200 ;
        RECT 0.985 71.760 131.000 75.800 ;
        RECT 4.400 70.360 131.000 71.760 ;
        RECT 0.985 66.320 131.000 70.360 ;
        RECT 4.400 64.920 131.000 66.320 ;
        RECT 0.985 63.600 131.000 64.920 ;
        RECT 0.985 62.200 130.600 63.600 ;
        RECT 0.985 60.880 131.000 62.200 ;
        RECT 4.400 59.480 131.000 60.880 ;
        RECT 0.985 55.440 131.000 59.480 ;
        RECT 4.400 54.040 131.000 55.440 ;
        RECT 0.985 50.000 131.000 54.040 ;
        RECT 4.400 48.600 131.000 50.000 ;
        RECT 0.985 45.920 131.000 48.600 ;
        RECT 0.985 44.560 130.600 45.920 ;
        RECT 4.400 44.520 130.600 44.560 ;
        RECT 4.400 43.160 131.000 44.520 ;
        RECT 0.985 39.120 131.000 43.160 ;
        RECT 4.400 37.720 131.000 39.120 ;
        RECT 0.985 33.680 131.000 37.720 ;
        RECT 4.400 32.280 131.000 33.680 ;
        RECT 0.985 28.240 131.000 32.280 ;
        RECT 4.400 26.840 130.600 28.240 ;
        RECT 0.985 22.800 131.000 26.840 ;
        RECT 4.400 21.400 131.000 22.800 ;
        RECT 0.985 17.360 131.000 21.400 ;
        RECT 4.400 15.960 131.000 17.360 ;
        RECT 0.985 11.920 131.000 15.960 ;
        RECT 4.400 10.560 131.000 11.920 ;
        RECT 4.400 10.520 130.600 10.560 ;
        RECT 0.985 9.160 130.600 10.520 ;
        RECT 0.985 6.480 131.000 9.160 ;
        RECT 4.400 5.275 131.000 6.480 ;
      LAYER met4 ;
        RECT 57.335 81.095 58.585 95.705 ;
  END
END dll
END LIBRARY

