VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO manual_routing
  CLASS COVER ;
  FOREIGN manual_routing ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.000 BY 1.000 ;
  PIN out
    PORT
      LAYER met2 ;
        RECT 1566.980 55.000 1568.255 56.270 ;
        RECT 1565.595 8.840 1569.595 55.000 ;
        RECT 1400.895 4.840 1569.595 8.840 ;
        RECT 1400.895 2.000 1404.895 4.840 ;
        RECT 1398.340 0.000 1407.320 2.000 ;
    END
    PORT
      LAYER met2 ;
        RECT 1466.980 55.000 1468.255 56.270 ;
        RECT 1465.610 15.620 1469.610 55.000 ;
        RECT 1290.870 11.620 1469.610 15.620 ;
        RECT 1290.870 2.000 1294.870 11.620 ;
        RECT 1288.340 0.000 1297.320 2.000 ;
    END
  END out
  PIN xi0_core
    PORT
      LAYER met2 ;
        RECT 944.945 29.030 948.915 30.020 ;
        RECT 944.930 15.530 948.930 29.030 ;
        RECT 944.930 11.530 1074.995 15.530 ;
        RECT 1070.995 2.000 1074.995 11.530 ;
        RECT 1068.340 0.000 1077.320 2.000 ;
      LAYER met3 ;
        RECT 946.555 30.000 947.315 31.295 ;
        RECT 944.965 28.070 948.895 30.000 ;
    END
  END xi0_core
  PIN xi1_core
    PORT
      LAYER met2 ;
        RECT 1288.340 0.000 1297.320 2.000 ;
    END
  END xi1_core
  PIN xo0_core
    PORT
      LAYER met2 ;
        RECT 1254.980 29.025 1258.950 30.020 ;
        RECT 1254.960 15.620 1258.960 29.025 ;
        RECT 1180.940 11.620 1258.960 15.620 ;
        RECT 1180.940 2.000 1184.940 11.620 ;
        RECT 1178.340 0.000 1187.320 2.000 ;
      LAYER met3 ;
        RECT 1256.555 30.000 1257.315 31.295 ;
        RECT 1255.000 28.070 1258.930 30.000 ;
    END
  END xo0_core
  PIN xo1_core
    PORT
      LAYER met2 ;
        RECT 1398.340 0.000 1407.320 2.000 ;
    END
  END xo1_core
  PIN adc_in
    PORT
      LAYER met3 ;
        RECT 1256.555 30.000 1257.315 31.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 946.555 30.000 947.315 31.265 ;
    END
  END adc_in
  PIN vssa3
    PORT
      LAYER met3 ;
        RECT 796.680 262.630 1700.260 272.630 ;
        RECT 1690.260 17.400 1700.260 262.630 ;
        RECT 1690.260 8.580 2365.645 17.400 ;
        RECT 1690.260 7.400 2365.655 8.580 ;
        RECT 2291.860 0.000 2315.760 7.400 ;
        RECT 2341.755 0.000 2365.655 7.400 ;
      LAYER met4 ;
        RECT 809.890 262.630 817.360 272.630 ;
        RECT 1119.890 262.630 1127.360 272.630 ;
        RECT 1495.850 211.255 1498.655 272.630 ;
        RECT 1595.850 211.255 1598.655 272.630 ;
        RECT 1649.430 159.560 1651.430 272.630 ;
      LAYER met5 ;
        RECT 809.890 232.235 817.360 272.630 ;
        RECT 1119.890 232.235 1127.360 272.630 ;
    END
  END vssa3
  PIN vdda3
    PORT
      LAYER met3 ;
        RECT 796.680 276.920 1713.400 286.920 ;
        RECT 1703.400 30.400 1713.400 276.920 ;
        RECT 1703.400 20.400 2495.655 30.400 ;
        RECT 2421.860 0.000 2445.760 20.400 ;
        RECT 2471.755 0.000 2495.655 20.400 ;
      LAYER met4 ;
        RECT 800.215 276.920 807.685 286.920 ;
        RECT 1110.215 276.920 1117.685 286.920 ;
        RECT 1499.510 211.255 1502.610 286.920 ;
        RECT 1599.510 211.255 1602.610 286.920 ;
        RECT 1652.980 159.560 1654.570 286.920 ;
      LAYER met5 ;
        RECT 800.215 232.235 807.685 286.920 ;
        RECT 1110.215 232.235 1117.685 286.920 ;
    END
  END vdda3
  PIN DVPWR
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1410.190 215.850 1426.495 217.760 ;
        RECT 1410.190 11.760 1412.100 215.850 ;
        RECT 1424.585 211.255 1426.495 215.850 ;
        RECT 1510.190 215.850 1526.495 217.760 ;
        RECT 1510.190 11.760 1512.100 215.850 ;
        RECT 1524.585 211.255 1526.495 215.850 ;
        RECT 1652.965 11.760 1654.610 100.005 ;
      LAYER met5 ;
        RECT 1085.460 19.760 1093.300 30.000 ;
        RECT 1395.460 19.760 1403.300 30.000 ;
        RECT 798.400 11.760 1688.800 19.760 ;
    END
  END DVPWR
  PIN DVGND
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1413.895 212.450 1419.910 214.360 ;
        RECT 1075.835 2.150 1083.675 37.840 ;
        RECT 1385.835 2.150 1393.675 37.840 ;
        RECT 1413.895 2.060 1415.805 212.450 ;
        RECT 1418.000 211.255 1419.910 212.450 ;
        RECT 1513.895 212.450 1519.910 214.360 ;
        RECT 1513.895 2.060 1515.805 212.450 ;
        RECT 1518.000 211.255 1519.910 212.450 ;
        RECT 1655.345 2.060 1656.575 100.005 ;
      LAYER met5 ;
        RECT 1075.835 30.000 1083.675 37.840 ;
        RECT 1385.835 30.000 1393.675 37.840 ;
        RECT 798.405 2.060 1688.800 10.060 ;
    END
  END DVGND
  OBS
      LAYER met2 ;
        RECT 798.725 273.905 1702.135 274.545 ;
        RECT 798.725 210.880 799.365 273.905 ;
        RECT 1108.760 210.880 1109.400 273.905 ;
        RECT 798.040 208.780 800.140 210.880 ;
        RECT 1108.040 208.780 1110.140 210.880 ;
        RECT 1701.495 19.245 1702.135 273.905 ;
        RECT 2661.895 47.140 2674.780 47.780 ;
        RECT 2661.895 19.245 2662.535 47.140 ;
        RECT 1701.495 18.605 2662.535 19.245 ;
      LAYER met3 ;
        RECT 798.040 208.780 800.140 210.880 ;
        RECT 1108.040 208.780 1110.140 210.880 ;
        RECT 1416.645 177.830 1418.205 178.830 ;
        RECT 1516.695 177.830 1518.255 178.830 ;
        RECT 1416.645 176.675 1417.645 177.830 ;
        RECT 1516.695 176.675 1517.695 177.830 ;
        RECT 1416.645 175.675 1418.220 176.675 ;
        RECT 1516.695 175.675 1518.270 176.675 ;
        RECT 1416.645 87.460 1418.205 88.460 ;
        RECT 1516.695 87.460 1518.255 88.460 ;
        RECT 1416.645 86.560 1417.645 87.460 ;
        RECT 1516.695 86.560 1517.695 87.460 ;
        RECT 1416.645 85.560 1418.220 86.560 ;
        RECT 1516.695 85.560 1518.270 86.560 ;
        RECT 812.120 30.750 814.900 31.745 ;
        RECT 1122.145 30.750 1124.925 31.745 ;
        RECT 812.120 30.110 878.405 30.750 ;
        RECT 1122.145 30.110 1188.430 30.750 ;
        RECT 812.120 28.965 814.900 30.110 ;
        RECT 1122.145 28.965 1124.925 30.110 ;
      LAYER met4 ;
        RECT 798.040 208.780 800.140 210.880 ;
        RECT 1108.040 208.780 1110.140 210.880 ;
        RECT 801.600 123.835 805.980 125.015 ;
        RECT 1111.560 123.835 1115.940 125.015 ;
        RECT 811.570 119.230 815.950 120.410 ;
        RECT 1121.530 119.230 1125.910 120.410 ;
        RECT 812.120 28.965 814.900 31.745 ;
        RECT 1122.145 28.965 1124.925 31.745 ;
      LAYER met5 ;
        RECT 801.480 123.625 806.100 125.225 ;
        RECT 1111.440 123.625 1116.060 125.225 ;
        RECT 811.450 119.020 816.070 120.620 ;
        RECT 1121.410 119.020 1126.030 120.620 ;
        RECT 812.000 28.845 815.020 31.865 ;
        RECT 1122.025 28.845 1125.045 31.865 ;
  END
END manual_routing
END LIBRARY

